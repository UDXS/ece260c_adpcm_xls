module adpcm_xls (clk,
    in_sample_rdy,
    in_sample_vld,
    out_pred_rdy,
    out_pred_vld,
    rst,
    in_sample,
    out_pred);
 input clk;
 output in_sample_rdy;
 input in_sample_vld;
 input out_pred_rdy;
 output out_pred_vld;
 input rst;
 input [15:0] in_sample;
 output [15:0] out_pred;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire clknet_0_clk;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0983_;
 wire _0985_;
 wire _0987_;
 wire _0989_;
 wire _0990_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1004_;
 wire _1009_;
 wire _1010_;
 wire _1012_;
 wire _1013_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire net239;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire net238;
 wire _1036_;
 wire _1037_;
 wire net237;
 wire net236;
 wire net235;
 wire net234;
 wire net233;
 wire net232;
 wire _1044_;
 wire net231;
 wire net230;
 wire net229;
 wire net228;
 wire _1049_;
 wire _1050_;
 wire net227;
 wire net226;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire net225;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire net223;
 wire net222;
 wire net221;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire net220;
 wire net219;
 wire net218;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire net217;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire net216;
 wire net215;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire net214;
 wire _1097_;
 wire _1098_;
 wire net213;
 wire _1100_;
 wire net212;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire net211;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire net210;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire net209;
 wire net208;
 wire net207;
 wire net206;
 wire _1178_;
 wire net205;
 wire net204;
 wire net203;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire net200;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire net188;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire net187;
 wire net186;
 wire net185;
 wire net184;
 wire net183;
 wire net182;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire net179;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire net178;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire net177;
 wire net176;
 wire net175;
 wire net174;
 wire net173;
 wire net172;
 wire _1560_;
 wire _1561_;
 wire net170;
 wire _1563_;
 wire _1564_;
 wire net168;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire clknet_3_1__leaf_clk;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire clknet_3_0__leaf_clk;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire net161;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire net160;
 wire _1676_;
 wire _1677_;
 wire net159;
 wire net158;
 wire net157;
 wire net156;
 wire net154;
 wire net153;
 wire net152;
 wire net151;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire net149;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire net148;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire net147;
 wire net146;
 wire net145;
 wire net144;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire net143;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire net135;
 wire net134;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire net133;
 wire net132;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire net129;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire net128;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire net125;
 wire _2001_;
 wire _2002_;
 wire net124;
 wire net123;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire net121;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire net120;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire net119;
 wire _2077_;
 wire net118;
 wire net117;
 wire net116;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire net115;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire net112;
 wire net111;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire net110;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire net109;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire net108;
 wire _2196_;
 wire net107;
 wire _2198_;
 wire net106;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire net104;
 wire net103;
 wire net102;
 wire net101;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire net100;
 wire net99;
 wire net98;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire net96;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire net95;
 wire _2230_;
 wire _2231_;
 wire net94;
 wire net93;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire net91;
 wire net90;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire net89;
 wire _2249_;
 wire _2250_;
 wire net88;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire net87;
 wire _2256_;
 wire _2257_;
 wire net86;
 wire net85;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire net81;
 wire _2298_;
 wire _2299_;
 wire net80;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire net78;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire net77;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire net74;
 wire net73;
 wire _2386_;
 wire net71;
 wire net70;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire net69;
 wire net68;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire net65;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire net64;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire net51;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire net50;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire net48;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire net47;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire net46;
 wire net45;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire net44;
 wire _2863_;
 wire _2864_;
 wire net43;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire net42;
 wire net41;
 wire net40;
 wire _2875_;
 wire _2876_;
 wire net39;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire net38;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire net37;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire net36;
 wire net35;
 wire net34;
 wire _2933_;
 wire net33;
 wire net32;
 wire net31;
 wire _2937_;
 wire net30;
 wire net29;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire net28;
 wire net27;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire net26;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire net25;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire net24;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire net23;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire net22;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire net21;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire net20;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire net19;
 wire _3081_;
 wire net18;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire net17;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire net16;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire net15;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire net166;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire net171;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire net181;
 wire _3205_;
 wire _3206_;
 wire net150;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire net192;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire net196;
 wire _3219_;
 wire net194;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire net131;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire net130;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire net201;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire net113;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire net76;
 wire net67;
 wire _3306_;
 wire net75;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire net62;
 wire _3312_;
 wire net61;
 wire _3314_;
 wire net97;
 wire _3316_;
 wire net84;
 wire _3318_;
 wire _3319_;
 wire net82;
 wire net57;
 wire _3322_;
 wire net55;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire net63;
 wire net105;
 wire net60;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire net92;
 wire net58;
 wire _3341_;
 wire net83;
 wire net56;
 wire _3344_;
 wire net79;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire net54;
 wire _3350_;
 wire net59;
 wire _3352_;
 wire net66;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire net224;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire net202;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire net199;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire net198;
 wire _3444_;
 wire net197;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire net195;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire net193;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire net191;
 wire _3470_;
 wire net190;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire net189;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire net180;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire net169;
 wire _3515_;
 wire net167;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire net165;
 wire _3522_;
 wire _3523_;
 wire net164;
 wire _3525_;
 wire net163;
 wire _3527_;
 wire _3528_;
 wire net162;
 wire _3530_;
 wire clknet_3_7__leaf_clk;
 wire _3532_;
 wire _3533_;
 wire clknet_3_6__leaf_clk;
 wire _3535_;
 wire clknet_3_5__leaf_clk;
 wire _3537_;
 wire _3538_;
 wire clknet_3_4__leaf_clk;
 wire _3540_;
 wire clknet_3_3__leaf_clk;
 wire _3542_;
 wire clknet_3_2__leaf_clk;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire net155;
 wire net142;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire net141;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire net140;
 wire _3591_;
 wire net139;
 wire _3593_;
 wire net138;
 wire _3595_;
 wire net137;
 wire net114;
 wire net136;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire net127;
 wire _3603_;
 wire net126;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire net122;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire net72;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire net52;
 wire net53;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire net49;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire \__in_sample_reg[10] ;
 wire \__in_sample_reg[11] ;
 wire \__in_sample_reg[12] ;
 wire \__in_sample_reg[13] ;
 wire \__in_sample_reg[14] ;
 wire \__in_sample_reg[15] ;
 wire \__in_sample_reg[1] ;
 wire \__in_sample_reg[2] ;
 wire \__in_sample_reg[3] ;
 wire \__in_sample_reg[4] ;
 wire \__in_sample_reg[5] ;
 wire \__in_sample_reg[6] ;
 wire \__in_sample_reg[7] ;
 wire \__in_sample_reg[8] ;
 wire \__in_sample_reg[9] ;
 wire \__st_0[0] ;
 wire \__st_0[10] ;
 wire \__st_0[11] ;
 wire \__st_0[12] ;
 wire \__st_0[13] ;
 wire \__st_0[1] ;
 wire \__st_0[2] ;
 wire \__st_0[3] ;
 wire \__st_0[4] ;
 wire \__st_0[6] ;
 wire \__st_0[7] ;
 wire \__st_0[8] ;
 wire \__st_0[9] ;
 wire \__st_1[0] ;
 wire \__st_1[10] ;
 wire \__st_1[11] ;
 wire \__st_1[12] ;
 wire \__st_1[13] ;
 wire \__st_1[14] ;
 wire \__st_1[15] ;
 wire \__st_1[16] ;
 wire \__st_1[17] ;
 wire \__st_1[18] ;
 wire \__st_1[19] ;
 wire \__st_1[20] ;
 wire \__st_1[21] ;
 wire \__st_1[22] ;
 wire \__st_1[23] ;
 wire \__st_1[24] ;
 wire \__st_1[25] ;
 wire \__st_1[26] ;
 wire \__st_1[27] ;
 wire \__st_1[28] ;
 wire \__st_1[29] ;
 wire \__st_1[2] ;
 wire \__st_1[3] ;
 wire \__st_1[4] ;
 wire \__st_1[5] ;
 wire \__st_1[6] ;
 wire \__st_1[7] ;
 wire \__st_1[8] ;
 wire \__st_1[9] ;
 wire \__st_2[0] ;
 wire \__st_2[10] ;
 wire \__st_2[11] ;
 wire \__st_2[12] ;
 wire \__st_2[13] ;
 wire \__st_2[1] ;
 wire \__st_2[2] ;
 wire \__st_2[3] ;
 wire \__st_2[4] ;
 wire \__st_2[6] ;
 wire \__st_2[7] ;
 wire \__st_2[8] ;
 wire \__st_2[9] ;
 wire net14;
 wire net6;
 wire net5;
 wire net4;
 wire net3;
 wire \__st_3[16] ;
 wire \__st_3[17] ;
 wire \__st_3[18] ;
 wire \__st_3[19] ;
 wire net13;
 wire \__st_3[20] ;
 wire \__st_3[21] ;
 wire \__st_3[22] ;
 wire \__st_3[23] ;
 wire \__st_3[24] ;
 wire \__st_3[25] ;
 wire \__st_3[26] ;
 wire \__st_3[27] ;
 wire \__st_3[28] ;
 wire \__st_3[29] ;
 wire net1;
 wire net2;
 wire net12;
 wire net11;
 wire net10;
 wire net9;
 wire net8;
 wire net7;

 INVx2_ASAP7_75t_R _3722_ (.A(_0546_),
    .Y(\__st_0[13] ));
 INVx2_ASAP7_75t_R _3723_ (.A(_3200_),
    .Y(\__st_0[12] ));
 INVx2_ASAP7_75t_R _3724_ (.A(_0547_),
    .Y(\__st_0[11] ));
 INVx2_ASAP7_75t_R _3725_ (.A(_3202_),
    .Y(\__st_0[10] ));
 INVx2_ASAP7_75t_R _3726_ (.A(_0548_),
    .Y(\__st_0[9] ));
 INVx2_ASAP7_75t_R _3727_ (.A(_0549_),
    .Y(\__st_0[8] ));
 INVx2_ASAP7_75t_R _3728_ (.A(_0550_),
    .Y(\__st_0[7] ));
 BUFx2_ASAP7_75t_R input12 (.A(in_sample[5]),
    .Y(net12));
 INVx2_ASAP7_75t_R _3730_ (.A(_0551_),
    .Y(\__st_0[6] ));
 INVx2_ASAP7_75t_R _3731_ (.A(_0553_),
    .Y(\__st_0[4] ));
 INVx2_ASAP7_75t_R _3732_ (.A(_0554_),
    .Y(\__st_0[3] ));
 INVx2_ASAP7_75t_R _3733_ (.A(_3206_),
    .Y(\__st_0[2] ));
 INVx2_ASAP7_75t_R _3734_ (.A(_0555_),
    .Y(\__st_0[1] ));
 BUFx2_ASAP7_75t_R input11 (.A(in_sample[4]),
    .Y(net11));
 INVx2_ASAP7_75t_R _3736_ (.A(_0556_),
    .Y(\__st_0[0] ));
 AND4x2_ASAP7_75t_R _3737_ (.A(_3202_),
    .B(_0548_),
    .C(_0549_),
    .D(_0550_),
    .Y(_0983_));
 BUFx2_ASAP7_75t_R input10 (.A(in_sample[3]),
    .Y(net10));
 AND4x2_ASAP7_75t_R _3739_ (.A(_3197_),
    .B(_0546_),
    .C(_3200_),
    .D(_0547_),
    .Y(_0985_));
 BUFx2_ASAP7_75t_R input9 (.A(in_sample[2]),
    .Y(net9));
 NAND2x2_ASAP7_75t_R _3741_ (.A(_0983_),
    .B(_0985_),
    .Y(_0987_));
 BUFx2_ASAP7_75t_R input8 (.A(in_sample[1]),
    .Y(net8));
 OR2x2_ASAP7_75t_R _3743_ (.A(\__st_0[6] ),
    .B(_0987_),
    .Y(_3403_));
 OR2x2_ASAP7_75t_R _3744_ (.A(_0553_),
    .B(_0554_),
    .Y(_0989_));
 AND3x2_ASAP7_75t_R _3745_ (.A(_3206_),
    .B(_0555_),
    .C(_0556_),
    .Y(_0990_));
 BUFx2_ASAP7_75t_R input7 (.A(in_sample[15]),
    .Y(net7));
 OA21x2_ASAP7_75t_R _3747_ (.A1(_0989_),
    .A2(_0990_),
    .B(_0552_),
    .Y(_0992_));
 AND2x2_ASAP7_75t_R _3748_ (.A(_0983_),
    .B(_0985_),
    .Y(_0993_));
 OA21x2_ASAP7_75t_R _3749_ (.A1(_0551_),
    .A2(_0992_),
    .B(_0993_),
    .Y(_0994_));
 INVx2_ASAP7_75t_R _3750_ (.A(_0994_),
    .Y(_0995_));
 OR2x2_ASAP7_75t_R _3751_ (.A(\__st_0[4] ),
    .B(_0995_),
    .Y(_3401_));
 AO21x2_ASAP7_75t_R _3752_ (.A1(\__st_0[2] ),
    .A2(_0994_),
    .B(_0243_),
    .Y(_0996_));
 OA21x2_ASAP7_75t_R _3753_ (.A1(\__st_0[3] ),
    .A2(_0995_),
    .B(_0996_),
    .Y(_3402_));
 OA21x2_ASAP7_75t_R _3754_ (.A1(_0553_),
    .A2(_0554_),
    .B(_0552_),
    .Y(_0997_));
 INVx2_ASAP7_75t_R _3755_ (.A(_0997_),
    .Y(_0998_));
 OA21x2_ASAP7_75t_R _3756_ (.A1(_0987_),
    .A2(_0998_),
    .B(_0996_),
    .Y(_0999_));
 INVx2_ASAP7_75t_R _3757_ (.A(_0552_),
    .Y(_1000_));
 AND4x2_ASAP7_75t_R _3758_ (.A(_0551_),
    .B(_1000_),
    .C(_0983_),
    .D(_0985_),
    .Y(_1001_));
 OR2x2_ASAP7_75t_R _3759_ (.A(_0999_),
    .B(_1001_),
    .Y(_3404_));
 BUFx2_ASAP7_75t_R input6 (.A(in_sample[14]),
    .Y(net6));
 BUFx2_ASAP7_75t_R input5 (.A(in_sample[13]),
    .Y(net5));
 XOR2x2_ASAP7_75t_R _3762_ (.A(_0698_),
    .B(_1001_),
    .Y(_1004_));
 BUFx2_ASAP7_75t_R input4 (.A(in_sample[12]),
    .Y(net4));
 BUFx2_ASAP7_75t_R input3 (.A(in_sample[11]),
    .Y(net3));
 TAPCELL_ASAP7_75t_R TAP_257 ();
 TAPCELL_ASAP7_75t_R TAP_256 ();
 INVx3_ASAP7_75t_R _3767_ (.A(_0697_),
    .Y(_1009_));
 OA21x2_ASAP7_75t_R _3768_ (.A1(_0551_),
    .A2(_0552_),
    .B(_0554_),
    .Y(_1010_));
 TAPCELL_ASAP7_75t_R TAP_255 ();
 AND3x2_ASAP7_75t_R _3770_ (.A(_0983_),
    .B(_0985_),
    .C(_1010_),
    .Y(_1012_));
 XNOR2x2_ASAP7_75t_R _3771_ (.A(_1009_),
    .B(_1012_),
    .Y(_1013_));
 TAPCELL_ASAP7_75t_R TAP_254 ();
 TAPCELL_ASAP7_75t_R TAP_253 ();
 TAPCELL_ASAP7_75t_R TAP_252 ();
 TAPCELL_ASAP7_75t_R TAP_251 ();
 TAPCELL_ASAP7_75t_R TAP_250 ();
 AND2x2_ASAP7_75t_R _3777_ (.A(net212),
    .B(net43),
    .Y(_1019_));
 AND2x2_ASAP7_75t_R _3778_ (.A(_1013_),
    .B(_1019_),
    .Y(_1020_));
 NAND2x2_ASAP7_75t_R _3779_ (.A(_1009_),
    .B(_1010_),
    .Y(_1021_));
 AO31x2_ASAP7_75t_R _3780_ (.A1(_0983_),
    .A2(_0985_),
    .A3(_1010_),
    .B(_1009_),
    .Y(_1022_));
 OA21x2_ASAP7_75t_R _3781_ (.A1(_0987_),
    .A2(_1021_),
    .B(_1022_),
    .Y(_1023_));
 CKINVDCx12_ASAP7_75t_R _3782_ (.A(net46),
    .Y(_1024_));
 CKINVDCx10_ASAP7_75t_R _3783_ (.A(net42),
    .Y(_1025_));
 TAPCELL_ASAP7_75t_R TAP_249 ();
 OR2x2_ASAP7_75t_R _3785_ (.A(_1024_),
    .B(_1025_),
    .Y(_1027_));
 AND2x2_ASAP7_75t_R _3786_ (.A(_1023_),
    .B(_1027_),
    .Y(_1028_));
 INVx2_ASAP7_75t_R _3787_ (.A(_0243_),
    .Y(_3399_));
 OA211x2_ASAP7_75t_R _3788_ (.A1(_0551_),
    .A2(_0997_),
    .B(_0985_),
    .C(_0983_),
    .Y(_1029_));
 OR2x6_ASAP7_75t_R _3789_ (.A(_3399_),
    .B(_1029_),
    .Y(_1030_));
 TAPCELL_ASAP7_75t_R TAP_248 ();
 OA21x2_ASAP7_75t_R _3791_ (.A1(_0551_),
    .A2(_0997_),
    .B(\__st_0[0] ),
    .Y(_1032_));
 AND2x6_ASAP7_75t_R _3792_ (.A(_0993_),
    .B(_1032_),
    .Y(_1033_));
 CKINVDCx10_ASAP7_75t_R _3793_ (.A(_1033_),
    .Y(_1034_));
 TAPCELL_ASAP7_75t_R TAP_247 ();
 AND2x2_ASAP7_75t_R _3795_ (.A(_1030_),
    .B(_1034_),
    .Y(_1036_));
 OA21x2_ASAP7_75t_R _3796_ (.A1(_1020_),
    .A2(_1028_),
    .B(_1036_),
    .Y(_1037_));
 TAPCELL_ASAP7_75t_R TAP_246 ();
 TAPCELL_ASAP7_75t_R TAP_245 ();
 TAPCELL_ASAP7_75t_R TAP_244 ();
 TAPCELL_ASAP7_75t_R TAP_243 ();
 TAPCELL_ASAP7_75t_R TAP_242 ();
 TAPCELL_ASAP7_75t_R TAP_241 ();
 OR2x2_ASAP7_75t_R _3803_ (.A(net43),
    .B(_1023_),
    .Y(_1044_));
 TAPCELL_ASAP7_75t_R TAP_240 ();
 TAPCELL_ASAP7_75t_R TAP_239 ();
 TAPCELL_ASAP7_75t_R TAP_238 ();
 TAPCELL_ASAP7_75t_R TAP_237 ();
 NOR2x2_ASAP7_75t_R _3808_ (.A(_0551_),
    .B(_0997_),
    .Y(_1049_));
 OA31x2_ASAP7_75t_R _3809_ (.A1(_0556_),
    .A2(_0987_),
    .A3(_1049_),
    .B1(net42),
    .Y(_1050_));
 TAPCELL_ASAP7_75t_R TAP_236 ();
 TAPCELL_ASAP7_75t_R TAP_235 ();
 OR2x2_ASAP7_75t_R _3812_ (.A(_1033_),
    .B(_1013_),
    .Y(_1053_));
 OA22x2_ASAP7_75t_R _3813_ (.A1(net46),
    .A2(_1050_),
    .B1(_1053_),
    .B2(_1027_),
    .Y(_1054_));
 OA21x2_ASAP7_75t_R _3814_ (.A1(_0987_),
    .A2(_1049_),
    .B(_0243_),
    .Y(_1055_));
 TAPCELL_ASAP7_75t_R TAP_234 ();
 AO21x2_ASAP7_75t_R _3816_ (.A1(_1044_),
    .A2(_1054_),
    .B(_1055_),
    .Y(_1057_));
 TAPCELL_ASAP7_75t_R TAP_233 ();
 AO21x2_ASAP7_75t_R _3818_ (.A1(net43),
    .A2(_1023_),
    .B(_1034_),
    .Y(_1058_));
 AO21x2_ASAP7_75t_R _3819_ (.A1(_1057_),
    .A2(_1058_),
    .B(net205),
    .Y(_1059_));
 INVx2_ASAP7_75t_R _3820_ (.A(_1059_),
    .Y(_1060_));
 AO21x2_ASAP7_75t_R _3821_ (.A1(net203),
    .A2(_1037_),
    .B(_1060_),
    .Y(_1061_));
 TAPCELL_ASAP7_75t_R TAP_232 ();
 TAPCELL_ASAP7_75t_R TAP_231 ();
 TAPCELL_ASAP7_75t_R TAP_230 ();
 AND2x2_ASAP7_75t_R _3825_ (.A(net43),
    .B(_1030_),
    .Y(_1065_));
 OA211x2_ASAP7_75t_R _3826_ (.A1(_1033_),
    .A2(_1065_),
    .B(_1023_),
    .C(net202),
    .Y(_1066_));
 AND2x2_ASAP7_75t_R _3827_ (.A(net199),
    .B(_1030_),
    .Y(_1067_));
 AND2x2_ASAP7_75t_R _3828_ (.A(_1033_),
    .B(_1023_),
    .Y(_1068_));
 AO21x2_ASAP7_75t_R _3829_ (.A1(_1013_),
    .A2(_1067_),
    .B(_1068_),
    .Y(_1069_));
 INVx13_ASAP7_75t_R _3830_ (.A(net41),
    .Y(_1070_));
 TAPCELL_ASAP7_75t_R TAP_229 ();
 TAPCELL_ASAP7_75t_R TAP_228 ();
 TAPCELL_ASAP7_75t_R TAP_227 ();
 AND2x2_ASAP7_75t_R _3834_ (.A(_1070_),
    .B(_1013_),
    .Y(_1074_));
 AND2x4_ASAP7_75t_R _3835_ (.A(_1025_),
    .B(_1033_),
    .Y(_1075_));
 AO221x2_ASAP7_75t_R _3836_ (.A1(net212),
    .A2(_1069_),
    .B1(_1074_),
    .B2(_1075_),
    .C(_1004_),
    .Y(_1076_));
 XNOR2x2_ASAP7_75t_R _3837_ (.A(_0698_),
    .B(_1001_),
    .Y(_1077_));
 OR3x2_ASAP7_75t_R _3838_ (.A(net197),
    .B(_1077_),
    .C(_1023_),
    .Y(_1078_));
 OR3x2_ASAP7_75t_R _3839_ (.A(_1033_),
    .B(_1065_),
    .C(_1078_),
    .Y(_1079_));
 INVx2_ASAP7_75t_R _3840_ (.A(_0459_),
    .Y(_1080_));
 OA211x2_ASAP7_75t_R _3841_ (.A1(_1066_),
    .A2(_1076_),
    .B(_1079_),
    .C(_1080_),
    .Y(_1081_));
 TAPCELL_ASAP7_75t_R TAP_226 ();
 AND2x2_ASAP7_75t_R _3843_ (.A(_1024_),
    .B(_1033_),
    .Y(_1083_));
 AO21x2_ASAP7_75t_R _3844_ (.A1(net43),
    .A2(_1070_),
    .B(_1013_),
    .Y(_1084_));
 AND2x2_ASAP7_75t_R _3845_ (.A(net43),
    .B(_1013_),
    .Y(_1085_));
 OA211x2_ASAP7_75t_R _3846_ (.A1(_0987_),
    .A2(_1021_),
    .B(_1022_),
    .C(_1025_),
    .Y(_1086_));
 OA21x2_ASAP7_75t_R _3847_ (.A1(_1070_),
    .A2(_1086_),
    .B(net215),
    .Y(_1087_));
 OA21x2_ASAP7_75t_R _3848_ (.A1(_1085_),
    .A2(_1087_),
    .B(_1034_),
    .Y(_1088_));
 AO21x2_ASAP7_75t_R _3849_ (.A1(_1083_),
    .A2(_1084_),
    .B(_1088_),
    .Y(_1089_));
 TAPCELL_ASAP7_75t_R TAP_225 ();
 TAPCELL_ASAP7_75t_R TAP_224 ();
 AO221x2_ASAP7_75t_R _3852_ (.A1(_1070_),
    .A2(_1013_),
    .B1(_1089_),
    .B2(_1030_),
    .C(_1077_),
    .Y(_1092_));
 AO32x2_ASAP7_75t_R _3853_ (.A1(_0459_),
    .A2(_1004_),
    .A3(_1061_),
    .B1(_1081_),
    .B2(_1092_),
    .Y(_1093_));
 NAND2x2_ASAP7_75t_R _3854_ (.A(_0700_),
    .B(_1093_),
    .Y(_3407_));
 INVx2_ASAP7_75t_R _3855_ (.A(_3407_),
    .Y(_3409_));
 AND2x4_ASAP7_75t_R _3856_ (.A(_1080_),
    .B(_0700_),
    .Y(_1094_));
 OA21x2_ASAP7_75t_R _3857_ (.A1(_3399_),
    .A2(_1029_),
    .B(net211),
    .Y(_1095_));
 TAPCELL_ASAP7_75t_R TAP_223 ();
 OA21x2_ASAP7_75t_R _3859_ (.A1(_1023_),
    .A2(_1050_),
    .B(_1095_),
    .Y(_1097_));
 OR2x4_ASAP7_75t_R _3860_ (.A(net41),
    .B(_1023_),
    .Y(_1098_));
 TAPCELL_ASAP7_75t_R TAP_222 ();
 OR4x2_ASAP7_75t_R _3862_ (.A(net43),
    .B(_0556_),
    .C(_0987_),
    .D(_1049_),
    .Y(_1100_));
 TAPCELL_ASAP7_75t_R TAP_221 ();
 OA21x2_ASAP7_75t_R _3864_ (.A1(net47),
    .A2(_1025_),
    .B(_1030_),
    .Y(_1102_));
 AND2x2_ASAP7_75t_R _3865_ (.A(_1100_),
    .B(_1102_),
    .Y(_1103_));
 AND2x2_ASAP7_75t_R _3866_ (.A(_0700_),
    .B(_1004_),
    .Y(_1104_));
 OA21x2_ASAP7_75t_R _3867_ (.A1(_1098_),
    .A2(_1103_),
    .B(_1104_),
    .Y(_1105_));
 INVx2_ASAP7_75t_R _3868_ (.A(_1050_),
    .Y(_1106_));
 OR2x2_ASAP7_75t_R _3869_ (.A(net41),
    .B(_1034_),
    .Y(_1107_));
 AO21x2_ASAP7_75t_R _3870_ (.A1(_1095_),
    .A2(_1107_),
    .B(net42),
    .Y(_1108_));
 AO21x2_ASAP7_75t_R _3871_ (.A1(_1106_),
    .A2(_1108_),
    .B(_1013_),
    .Y(_1109_));
 OA211x2_ASAP7_75t_R _3872_ (.A1(_1070_),
    .A2(_1097_),
    .B(_1105_),
    .C(_1109_),
    .Y(_1110_));
 AO21x2_ASAP7_75t_R _3873_ (.A1(_1030_),
    .A2(_1027_),
    .B(_1033_),
    .Y(_1111_));
 AND2x2_ASAP7_75t_R _3874_ (.A(_1100_),
    .B(_1111_),
    .Y(_1112_));
 TAPCELL_ASAP7_75t_R TAP_220 ();
 OR2x2_ASAP7_75t_R _3876_ (.A(_1025_),
    .B(_1023_),
    .Y(_1114_));
 OR2x2_ASAP7_75t_R _3877_ (.A(net42),
    .B(_1070_),
    .Y(_1115_));
 AO21x2_ASAP7_75t_R _3878_ (.A1(net47),
    .A2(_1013_),
    .B(_1115_),
    .Y(_1116_));
 OA21x2_ASAP7_75t_R _3879_ (.A1(_1024_),
    .A2(_1114_),
    .B(_1116_),
    .Y(_1117_));
 AO21x2_ASAP7_75t_R _3880_ (.A1(_1034_),
    .A2(_1013_),
    .B(net47),
    .Y(_1118_));
 AO21x2_ASAP7_75t_R _3881_ (.A1(net41),
    .A2(_1118_),
    .B(_1025_),
    .Y(_1119_));
 OA21x2_ASAP7_75t_R _3882_ (.A1(_1033_),
    .A2(_1117_),
    .B(_1119_),
    .Y(_1120_));
 AND2x2_ASAP7_75t_R _3883_ (.A(_1034_),
    .B(_1023_),
    .Y(_1121_));
 NOR2x2_ASAP7_75t_R _3884_ (.A(_0697_),
    .B(_1010_),
    .Y(_1122_));
 AND2x2_ASAP7_75t_R _3885_ (.A(_0697_),
    .B(_1010_),
    .Y(_1123_));
 OR5x2_ASAP7_75t_R _3886_ (.A(_0556_),
    .B(_0987_),
    .C(_1049_),
    .D(_1122_),
    .E(_1123_),
    .Y(_1124_));
 OA22x2_ASAP7_75t_R _3887_ (.A1(net200),
    .A2(_1121_),
    .B1(_1124_),
    .B2(net43),
    .Y(_1125_));
 OA21x2_ASAP7_75t_R _3888_ (.A1(_1055_),
    .A2(_1120_),
    .B(_1125_),
    .Y(_1126_));
 INVx2_ASAP7_75t_R _3889_ (.A(_1126_),
    .Y(_1127_));
 OA211x2_ASAP7_75t_R _3890_ (.A1(_1098_),
    .A2(_1112_),
    .B(_1127_),
    .C(_1004_),
    .Y(_1128_));
 OR2x2_ASAP7_75t_R _3891_ (.A(_1034_),
    .B(_1013_),
    .Y(_1129_));
 OA21x2_ASAP7_75t_R _3892_ (.A1(net42),
    .A2(_1023_),
    .B(_1129_),
    .Y(_1130_));
 OA21x2_ASAP7_75t_R _3893_ (.A1(net46),
    .A2(_1130_),
    .B(_1112_),
    .Y(_1131_));
 OR2x6_ASAP7_75t_R _3894_ (.A(net41),
    .B(_1013_),
    .Y(_1132_));
 TAPCELL_ASAP7_75t_R TAP_219 ();
 AND2x2_ASAP7_75t_R _3896_ (.A(_1024_),
    .B(_1030_),
    .Y(_1134_));
 OR2x2_ASAP7_75t_R _3897_ (.A(net46),
    .B(net42),
    .Y(_1135_));
 OA21x2_ASAP7_75t_R _3898_ (.A1(_1033_),
    .A2(_1134_),
    .B(_1135_),
    .Y(_1136_));
 OA21x2_ASAP7_75t_R _3899_ (.A1(_1132_),
    .A2(_1136_),
    .B(_1077_),
    .Y(_1137_));
 AND2x2_ASAP7_75t_R _3900_ (.A(net43),
    .B(_1033_),
    .Y(_1138_));
 AO21x2_ASAP7_75t_R _3901_ (.A1(_1025_),
    .A2(_1036_),
    .B(_1138_),
    .Y(_1139_));
 OR2x2_ASAP7_75t_R _3902_ (.A(_1050_),
    .B(_1075_),
    .Y(_1140_));
 AO221x2_ASAP7_75t_R _3903_ (.A1(net210),
    .A2(_1139_),
    .B1(_1134_),
    .B2(_1140_),
    .C(_1098_),
    .Y(_1141_));
 OA211x2_ASAP7_75t_R _3904_ (.A1(_1070_),
    .A2(_1131_),
    .B(_1137_),
    .C(_1141_),
    .Y(_1142_));
 OR3x2_ASAP7_75t_R _3905_ (.A(_0459_),
    .B(_1128_),
    .C(_1142_),
    .Y(_1143_));
 OA21x2_ASAP7_75t_R _3906_ (.A1(_1094_),
    .A2(_1110_),
    .B(_1143_),
    .Y(_3217_));
 INVx2_ASAP7_75t_R _3907_ (.A(_3217_),
    .Y(_3174_));
 CKINVDCx14_ASAP7_75t_R _3908_ (.A(_3145_),
    .Y(\__in_sample_reg[15] ));
 OA21x2_ASAP7_75t_R _3909_ (.A1(_0451_),
    .A2(_0452_),
    .B(_0450_),
    .Y(_1144_));
 OA21x2_ASAP7_75t_R _3910_ (.A1(_0706_),
    .A2(_1144_),
    .B(_0449_),
    .Y(_3130_));
 OA21x2_ASAP7_75t_R _3911_ (.A1(_0448_),
    .A2(_3130_),
    .B(_0447_),
    .Y(_1145_));
 OA21x2_ASAP7_75t_R _3912_ (.A1(_0446_),
    .A2(_1145_),
    .B(_0445_),
    .Y(_1146_));
 OA21x2_ASAP7_75t_R _3913_ (.A1(_0444_),
    .A2(_1146_),
    .B(_0443_),
    .Y(_1147_));
 OA21x2_ASAP7_75t_R _3914_ (.A1(_0705_),
    .A2(_1147_),
    .B(_0442_),
    .Y(_1148_));
 OA21x2_ASAP7_75t_R _3915_ (.A1(_0441_),
    .A2(_1148_),
    .B(_0440_),
    .Y(_1149_));
 AND3x2_ASAP7_75t_R _3916_ (.A(_0437_),
    .B(_0436_),
    .C(_0439_),
    .Y(_1150_));
 OA21x2_ASAP7_75t_R _3917_ (.A1(_0704_),
    .A2(_1149_),
    .B(_1150_),
    .Y(_1151_));
 AND3x2_ASAP7_75t_R _3918_ (.A(_0437_),
    .B(_0436_),
    .C(_0438_),
    .Y(_1152_));
 AO21x2_ASAP7_75t_R _3919_ (.A1(_0436_),
    .A2(_0703_),
    .B(_1152_),
    .Y(_1153_));
 OR3x2_ASAP7_75t_R _3920_ (.A(_0432_),
    .B(_0435_),
    .C(_0702_),
    .Y(_1154_));
 OR3x2_ASAP7_75t_R _3921_ (.A(_0432_),
    .B(_0434_),
    .C(_0702_),
    .Y(_1155_));
 OA21x2_ASAP7_75t_R _3922_ (.A1(_0432_),
    .A2(_0433_),
    .B(_1155_),
    .Y(_1156_));
 OA31x2_ASAP7_75t_R _3923_ (.A1(_1151_),
    .A2(_1153_),
    .A3(_1154_),
    .B1(_1156_),
    .Y(_1157_));
 AND2x2_ASAP7_75t_R _3924_ (.A(_0431_),
    .B(_1157_),
    .Y(_1158_));
 OA21x2_ASAP7_75t_R _3925_ (.A1(net173),
    .A2(_1158_),
    .B(_0429_),
    .Y(_3150_));
 AND3x2_ASAP7_75t_R _3926_ (.A(_0426_),
    .B(_0424_),
    .C(_0429_),
    .Y(_1159_));
 OA21x2_ASAP7_75t_R _3927_ (.A1(_0422_),
    .A2(_0421_),
    .B(_0420_),
    .Y(_1160_));
 AND3x2_ASAP7_75t_R _3928_ (.A(_0431_),
    .B(_1159_),
    .C(_1160_),
    .Y(_1161_));
 AO21x2_ASAP7_75t_R _3929_ (.A1(_0430_),
    .A2(_0429_),
    .B(_0428_),
    .Y(_1162_));
 AO21x2_ASAP7_75t_R _3930_ (.A1(_0426_),
    .A2(_1162_),
    .B(_0425_),
    .Y(_1163_));
 AND2x2_ASAP7_75t_R _3931_ (.A(_0424_),
    .B(_1163_),
    .Y(_1164_));
 OR3x2_ASAP7_75t_R _3932_ (.A(_0421_),
    .B(_0423_),
    .C(_1164_),
    .Y(_1165_));
 AO21x2_ASAP7_75t_R _3933_ (.A1(_1160_),
    .A2(_1165_),
    .B(_0419_),
    .Y(_1166_));
 AO21x2_ASAP7_75t_R _3934_ (.A1(_1157_),
    .A2(_1161_),
    .B(_1166_),
    .Y(_1167_));
 AND3x2_ASAP7_75t_R _3935_ (.A(_0413_),
    .B(_0418_),
    .C(_0416_),
    .Y(_1168_));
 AND3x2_ASAP7_75t_R _3936_ (.A(_0413_),
    .B(_0417_),
    .C(_0416_),
    .Y(_1169_));
 AO221x2_ASAP7_75t_R _3937_ (.A1(_0413_),
    .A2(_0415_),
    .B1(_1167_),
    .B2(_1168_),
    .C(_1169_),
    .Y(_1170_));
 OA21x2_ASAP7_75t_R _3938_ (.A1(_0410_),
    .A2(_1170_),
    .B(_0409_),
    .Y(_3146_));
 INVx2_ASAP7_75t_R _3939_ (.A(_0567_),
    .Y(_1171_));
 XNOR2x2_ASAP7_75t_R _3940_ (.A(_0453_),
    .B(_3145_),
    .Y(_1172_));
 XNOR2x2_ASAP7_75t_R _3941_ (.A(_1171_),
    .B(_1172_),
    .Y(_1173_));
 TAPCELL_ASAP7_75t_R TAP_218 ();
 TAPCELL_ASAP7_75t_R TAP_217 ();
 TAPCELL_ASAP7_75t_R TAP_216 ();
 TAPCELL_ASAP7_75t_R TAP_215 ();
 XNOR2x2_ASAP7_75t_R _3946_ (.A(_0567_),
    .B(_1172_),
    .Y(_1178_));
 TAPCELL_ASAP7_75t_R TAP_214 ();
 TAPCELL_ASAP7_75t_R TAP_213 ();
 TAPCELL_ASAP7_75t_R TAP_212 ();
 AND2x2_ASAP7_75t_R _3950_ (.A(_0454_),
    .B(net227),
    .Y(_1182_));
 AO21x2_ASAP7_75t_R _3951_ (.A1(_3427_),
    .A2(_1173_),
    .B(_1182_),
    .Y(_1183_));
 TAPCELL_ASAP7_75t_R TAP_211 ();
 OR2x2_ASAP7_75t_R _3953_ (.A(_1024_),
    .B(_1033_),
    .Y(_1184_));
 AO21x2_ASAP7_75t_R _3954_ (.A1(_1065_),
    .A2(_1184_),
    .B(_1098_),
    .Y(_1185_));
 AO21x2_ASAP7_75t_R _3955_ (.A1(_1023_),
    .A2(_1111_),
    .B(_1070_),
    .Y(_1186_));
 OR2x2_ASAP7_75t_R _3956_ (.A(_1024_),
    .B(net43),
    .Y(_1187_));
 AO221x2_ASAP7_75t_R _3957_ (.A1(net46),
    .A2(_1075_),
    .B1(_1187_),
    .B2(_1036_),
    .C(_1132_),
    .Y(_1188_));
 AND4x2_ASAP7_75t_R _3958_ (.A(_1104_),
    .B(_1185_),
    .C(_1186_),
    .D(_1188_),
    .Y(_1189_));
 AND2x2_ASAP7_75t_R _3959_ (.A(net42),
    .B(net41),
    .Y(_1190_));
 AO221x2_ASAP7_75t_R _3960_ (.A1(_1025_),
    .A2(_1034_),
    .B1(_1190_),
    .B2(net47),
    .C(_1023_),
    .Y(_1191_));
 OA21x2_ASAP7_75t_R _3961_ (.A1(net47),
    .A2(_1050_),
    .B(_1023_),
    .Y(_1192_));
 INVx2_ASAP7_75t_R _3962_ (.A(_1192_),
    .Y(_1193_));
 AND4x2_ASAP7_75t_R _3963_ (.A(_1077_),
    .B(_1030_),
    .C(_1191_),
    .D(_1193_),
    .Y(_1194_));
 AND2x2_ASAP7_75t_R _3964_ (.A(_1034_),
    .B(_1095_),
    .Y(_1195_));
 OR3x2_ASAP7_75t_R _3965_ (.A(_1065_),
    .B(_1098_),
    .C(_1195_),
    .Y(_1196_));
 OR2x2_ASAP7_75t_R _3966_ (.A(_1024_),
    .B(_1034_),
    .Y(_1197_));
 AO221x2_ASAP7_75t_R _3967_ (.A1(net212),
    .A2(_1075_),
    .B1(_1197_),
    .B2(_1065_),
    .C(_1132_),
    .Y(_1198_));
 OA21x2_ASAP7_75t_R _3968_ (.A1(_1033_),
    .A2(_1023_),
    .B(_1025_),
    .Y(_1199_));
 OA211x2_ASAP7_75t_R _3969_ (.A1(net46),
    .A2(_1053_),
    .B(_1124_),
    .C(net43),
    .Y(_1200_));
 OA21x2_ASAP7_75t_R _3970_ (.A1(_1024_),
    .A2(_1050_),
    .B(_1030_),
    .Y(_1201_));
 OA21x2_ASAP7_75t_R _3971_ (.A1(_1199_),
    .A2(_1200_),
    .B(_1201_),
    .Y(_1202_));
 AND2x2_ASAP7_75t_R _3972_ (.A(_1033_),
    .B(_1086_),
    .Y(_1203_));
 OR3x2_ASAP7_75t_R _3973_ (.A(_1070_),
    .B(_1202_),
    .C(_1203_),
    .Y(_1204_));
 AND4x2_ASAP7_75t_R _3974_ (.A(_1004_),
    .B(_1196_),
    .C(_1198_),
    .D(_1204_),
    .Y(_1205_));
 OR3x2_ASAP7_75t_R _3975_ (.A(_0459_),
    .B(_1194_),
    .C(_1205_),
    .Y(_1206_));
 OA21x2_ASAP7_75t_R _3976_ (.A1(_1094_),
    .A2(_1189_),
    .B(_1206_),
    .Y(_1207_));
 TAPCELL_ASAP7_75t_R TAP_210 ();
 INVx3_ASAP7_75t_R _3978_ (.A(_1207_),
    .Y(_3180_));
 XNOR2x2_ASAP7_75t_R _3979_ (.A(_0455_),
    .B(_0706_),
    .Y(_1208_));
 TAPCELL_ASAP7_75t_R TAP_209 ();
 AND2x2_ASAP7_75t_R _3981_ (.A(_0456_),
    .B(net239),
    .Y(_1210_));
 XOR2x2_ASAP7_75t_R _3982_ (.A(_1208_),
    .B(_1210_),
    .Y(_3430_));
 OR2x2_ASAP7_75t_R _3983_ (.A(_1075_),
    .B(_1132_),
    .Y(_1211_));
 AO21x2_ASAP7_75t_R _3984_ (.A1(net43),
    .A2(_1134_),
    .B(_1211_),
    .Y(_1212_));
 OA21x2_ASAP7_75t_R _3985_ (.A1(_3399_),
    .A2(_1029_),
    .B(_1025_),
    .Y(_1213_));
 OA21x2_ASAP7_75t_R _3986_ (.A1(_1138_),
    .A2(_1213_),
    .B(net218),
    .Y(_1214_));
 AND2x2_ASAP7_75t_R _3987_ (.A(_1024_),
    .B(net42),
    .Y(_1215_));
 AO21x2_ASAP7_75t_R _3988_ (.A1(_1036_),
    .A2(_1215_),
    .B(_1098_),
    .Y(_1216_));
 OA211x2_ASAP7_75t_R _3989_ (.A1(_1214_),
    .A2(_1216_),
    .B(_0459_),
    .C(_1004_),
    .Y(_1217_));
 XNOR2x2_ASAP7_75t_R _3990_ (.A(_1023_),
    .B(_1184_),
    .Y(_1218_));
 AO21x2_ASAP7_75t_R _3991_ (.A1(_1065_),
    .A2(_1218_),
    .B(_1070_),
    .Y(_1219_));
 AND3x2_ASAP7_75t_R _3992_ (.A(_1036_),
    .B(_1013_),
    .C(_1135_),
    .Y(_1220_));
 OA211x2_ASAP7_75t_R _3993_ (.A1(_1033_),
    .A2(_1095_),
    .B(net42),
    .C(net41),
    .Y(_1221_));
 AO21x2_ASAP7_75t_R _3994_ (.A1(_1070_),
    .A2(_1220_),
    .B(_1221_),
    .Y(_1222_));
 OA31x2_ASAP7_75t_R _3995_ (.A1(_0556_),
    .A2(_0987_),
    .A3(_1049_),
    .B1(_1025_),
    .Y(_1223_));
 OA21x2_ASAP7_75t_R _3996_ (.A1(_1024_),
    .A2(_1223_),
    .B(_1030_),
    .Y(_1224_));
 OR4x2_ASAP7_75t_R _3997_ (.A(_1025_),
    .B(net41),
    .C(_1033_),
    .D(_1220_),
    .Y(_1225_));
 OA21x2_ASAP7_75t_R _3998_ (.A1(_1013_),
    .A2(_1224_),
    .B(_1225_),
    .Y(_1226_));
 OA21x2_ASAP7_75t_R _3999_ (.A1(_1023_),
    .A2(_1222_),
    .B(_1226_),
    .Y(_1227_));
 AO21x2_ASAP7_75t_R _4000_ (.A1(_1030_),
    .A2(_1135_),
    .B(_1070_),
    .Y(_1228_));
 INVx2_ASAP7_75t_R _4001_ (.A(_1107_),
    .Y(_1229_));
 AO21x2_ASAP7_75t_R _4002_ (.A1(net42),
    .A2(_1229_),
    .B(_1223_),
    .Y(_1230_));
 AO32x2_ASAP7_75t_R _4003_ (.A1(net42),
    .A2(_1034_),
    .A3(_1098_),
    .B1(_1230_),
    .B2(_1024_),
    .Y(_1231_));
 OA21x2_ASAP7_75t_R _4004_ (.A1(net47),
    .A2(_1013_),
    .B(_1229_),
    .Y(_1232_));
 AO222x2_ASAP7_75t_R _4005_ (.A1(net41),
    .A2(_1023_),
    .B1(_1231_),
    .B2(_1030_),
    .C1(_1232_),
    .C2(_1025_),
    .Y(_1233_));
 OA211x2_ASAP7_75t_R _4006_ (.A1(_1053_),
    .A2(_1228_),
    .B(_1233_),
    .C(_1004_),
    .Y(_1234_));
 AO21x2_ASAP7_75t_R _4007_ (.A1(_1077_),
    .A2(_1227_),
    .B(_1234_),
    .Y(_1235_));
 AO32x2_ASAP7_75t_R _4008_ (.A1(_1212_),
    .A2(_1217_),
    .A3(_1219_),
    .B1(_1235_),
    .B2(_1080_),
    .Y(_1236_));
 AND2x6_ASAP7_75t_R _4009_ (.A(_0700_),
    .B(_1236_),
    .Y(_3233_));
 INVx4_ASAP7_75t_R _4010_ (.A(_3233_),
    .Y(_3171_));
 AND2x2_ASAP7_75t_R _4011_ (.A(_0457_),
    .B(net227),
    .Y(_1237_));
 AO21x2_ASAP7_75t_R _4012_ (.A1(_3433_),
    .A2(_1173_),
    .B(_1237_),
    .Y(_1238_));
 TAPCELL_ASAP7_75t_R TAP_208 ();
 AND2x2_ASAP7_75t_R _4014_ (.A(_1004_),
    .B(_1094_),
    .Y(_1239_));
 AND3x2_ASAP7_75t_R _4015_ (.A(_1024_),
    .B(_1033_),
    .C(_1023_),
    .Y(_1240_));
 OA211x2_ASAP7_75t_R _4016_ (.A1(net212),
    .A2(_1034_),
    .B(_1013_),
    .C(_1030_),
    .Y(_1241_));
 OA21x2_ASAP7_75t_R _4017_ (.A1(_1240_),
    .A2(_1241_),
    .B(_0263_),
    .Y(_1242_));
 AO21x2_ASAP7_75t_R _4018_ (.A1(_1023_),
    .A2(_1213_),
    .B(_1070_),
    .Y(_1243_));
 OA211x2_ASAP7_75t_R _4019_ (.A1(net47),
    .A2(_1223_),
    .B(_1013_),
    .C(_1030_),
    .Y(_1244_));
 AND3x2_ASAP7_75t_R _4020_ (.A(_0993_),
    .B(_1032_),
    .C(_1135_),
    .Y(_1245_));
 AO21x2_ASAP7_75t_R _4021_ (.A1(_1023_),
    .A2(_1245_),
    .B(net198),
    .Y(_1246_));
 OA21x2_ASAP7_75t_R _4022_ (.A1(_1244_),
    .A2(_1246_),
    .B(_1094_),
    .Y(_1247_));
 OA21x2_ASAP7_75t_R _4023_ (.A1(_1242_),
    .A2(_1243_),
    .B(_1247_),
    .Y(_1248_));
 OR3x2_ASAP7_75t_R _4024_ (.A(net46),
    .B(_1033_),
    .C(_1023_),
    .Y(_1249_));
 AO21x2_ASAP7_75t_R _4025_ (.A1(_1129_),
    .A2(_1249_),
    .B(_1025_),
    .Y(_1250_));
 OA21x2_ASAP7_75t_R _4026_ (.A1(_3399_),
    .A2(_1029_),
    .B(_1070_),
    .Y(_1251_));
 OA211x2_ASAP7_75t_R _4027_ (.A1(net43),
    .A2(_1053_),
    .B(_1197_),
    .C(_1251_),
    .Y(_1252_));
 AND2x2_ASAP7_75t_R _4028_ (.A(_1024_),
    .B(_1025_),
    .Y(_1253_));
 XNOR2x2_ASAP7_75t_R _4029_ (.A(_1024_),
    .B(_1033_),
    .Y(_1254_));
 OR2x2_ASAP7_75t_R _4030_ (.A(net43),
    .B(_1013_),
    .Y(_1255_));
 AO221x2_ASAP7_75t_R _4031_ (.A1(_1121_),
    .A2(_1253_),
    .B1(_1254_),
    .B2(_1255_),
    .C(_1085_),
    .Y(_1256_));
 AO221x2_ASAP7_75t_R _4032_ (.A1(_1250_),
    .A2(_1252_),
    .B1(_1256_),
    .B2(_1067_),
    .C(_1077_),
    .Y(_1257_));
 OA21x2_ASAP7_75t_R _4033_ (.A1(_1239_),
    .A2(_1248_),
    .B(_1257_),
    .Y(_3436_));
 INVx5_ASAP7_75t_R _4034_ (.A(_3436_),
    .Y(_3182_));
 INVx2_ASAP7_75t_R _4035_ (.A(_0707_),
    .Y(_3428_));
 AND3x2_ASAP7_75t_R _4036_ (.A(_3433_),
    .B(_3428_),
    .C(_1208_),
    .Y(_3450_));
 XOR2x2_ASAP7_75t_R _4037_ (.A(_0446_),
    .B(_0461_),
    .Y(_1258_));
 AND3x2_ASAP7_75t_R _4038_ (.A(_3449_),
    .B(_3450_),
    .C(_1258_),
    .Y(_3441_));
 XNOR2x2_ASAP7_75t_R _4039_ (.A(_0460_),
    .B(_0705_),
    .Y(_1259_));
 AND2x2_ASAP7_75t_R _4040_ (.A(_0462_),
    .B(net239),
    .Y(_1260_));
 XOR2x2_ASAP7_75t_R _4041_ (.A(_1259_),
    .B(_1260_),
    .Y(_3437_));
 OR3x2_ASAP7_75t_R _4042_ (.A(net216),
    .B(_0556_),
    .C(_1049_),
    .Y(_1261_));
 AND4x2_ASAP7_75t_R _4043_ (.A(_0697_),
    .B(_0983_),
    .C(_0985_),
    .D(_1010_),
    .Y(_1262_));
 OR2x2_ASAP7_75t_R _4044_ (.A(_1262_),
    .B(_1122_),
    .Y(_1263_));
 AND2x2_ASAP7_75t_R _4045_ (.A(_1009_),
    .B(_0987_),
    .Y(_1264_));
 AO221x2_ASAP7_75t_R _4046_ (.A1(net216),
    .A2(_1223_),
    .B1(_1261_),
    .B2(_1263_),
    .C(_1264_),
    .Y(_1265_));
 AND2x2_ASAP7_75t_R _4047_ (.A(_1013_),
    .B(_1215_),
    .Y(_1266_));
 OA21x2_ASAP7_75t_R _4048_ (.A1(_1265_),
    .A2(_1266_),
    .B(_1030_),
    .Y(_1267_));
 AO21x2_ASAP7_75t_R _4049_ (.A1(_1013_),
    .A2(_1138_),
    .B(net199),
    .Y(_1268_));
 AO21x2_ASAP7_75t_R _4050_ (.A1(_1053_),
    .A2(_1124_),
    .B(_1115_),
    .Y(_1269_));
 OR2x2_ASAP7_75t_R _4051_ (.A(_1070_),
    .B(_1033_),
    .Y(_1270_));
 OA21x2_ASAP7_75t_R _4052_ (.A1(_1102_),
    .A2(_1270_),
    .B(_1004_),
    .Y(_1271_));
 OA211x2_ASAP7_75t_R _4053_ (.A1(_1267_),
    .A2(_1268_),
    .B(_1269_),
    .C(_1271_),
    .Y(_1272_));
 AND2x2_ASAP7_75t_R _4054_ (.A(_1033_),
    .B(_1190_),
    .Y(_1273_));
 AND2x2_ASAP7_75t_R _4055_ (.A(_1025_),
    .B(_1070_),
    .Y(_1274_));
 AND3x2_ASAP7_75t_R _4056_ (.A(_1034_),
    .B(_1023_),
    .C(_1274_),
    .Y(_1275_));
 OA211x2_ASAP7_75t_R _4057_ (.A1(_1273_),
    .A2(_1275_),
    .B(_1077_),
    .C(_1134_),
    .Y(_1276_));
 AO21x2_ASAP7_75t_R _4058_ (.A1(_1009_),
    .A2(_0987_),
    .B(_1262_),
    .Y(_1277_));
 NAND2x2_ASAP7_75t_R _4059_ (.A(_1024_),
    .B(_1277_),
    .Y(_1278_));
 AND2x2_ASAP7_75t_R _4060_ (.A(_1024_),
    .B(_1190_),
    .Y(_1279_));
 OR3x2_ASAP7_75t_R _4061_ (.A(net210),
    .B(_0697_),
    .C(_1010_),
    .Y(_1280_));
 OA211x2_ASAP7_75t_R _4062_ (.A1(_1274_),
    .A2(_1279_),
    .B(_1280_),
    .C(_1033_),
    .Y(_1281_));
 AND3x2_ASAP7_75t_R _4063_ (.A(_1077_),
    .B(_1278_),
    .C(_1281_),
    .Y(_1282_));
 OR3x2_ASAP7_75t_R _4064_ (.A(_1025_),
    .B(_1070_),
    .C(_1023_),
    .Y(_1283_));
 OR4x2_ASAP7_75t_R _4065_ (.A(_1025_),
    .B(_0556_),
    .C(_0987_),
    .D(_1049_),
    .Y(_1284_));
 AND3x2_ASAP7_75t_R _4066_ (.A(_1077_),
    .B(_1030_),
    .C(_1284_),
    .Y(_1285_));
 OR2x2_ASAP7_75t_R _4067_ (.A(net42),
    .B(net41),
    .Y(_1286_));
 AO21x2_ASAP7_75t_R _4068_ (.A1(_1013_),
    .A2(_1286_),
    .B(net47),
    .Y(_1287_));
 AND4x2_ASAP7_75t_R _4069_ (.A(_1132_),
    .B(_1283_),
    .C(_1285_),
    .D(_1287_),
    .Y(_1288_));
 OR4x2_ASAP7_75t_R _4070_ (.A(_0459_),
    .B(_1276_),
    .C(_1282_),
    .D(_1288_),
    .Y(_1289_));
 AND4x2_ASAP7_75t_R _4071_ (.A(_1070_),
    .B(_0700_),
    .C(_1004_),
    .D(_1095_),
    .Y(_1290_));
 AO32x2_ASAP7_75t_R _4072_ (.A1(net43),
    .A2(_1023_),
    .A3(_1290_),
    .B1(_1080_),
    .B2(_0700_),
    .Y(_1291_));
 OA21x2_ASAP7_75t_R _4073_ (.A1(_1272_),
    .A2(_1289_),
    .B(_1291_),
    .Y(_3442_));
 INVx4_ASAP7_75t_R _4074_ (.A(_3442_),
    .Y(_3165_));
 AND2x2_ASAP7_75t_R _4075_ (.A(_0463_),
    .B(net237),
    .Y(_1292_));
 AO21x2_ASAP7_75t_R _4076_ (.A1(_3440_),
    .A2(_1173_),
    .B(_1292_),
    .Y(_1293_));
 TAPCELL_ASAP7_75t_R TAP_207 ();
 AND3x2_ASAP7_75t_R _4078_ (.A(_1034_),
    .B(_1013_),
    .C(_1019_),
    .Y(_1294_));
 AND2x2_ASAP7_75t_R _4079_ (.A(_0459_),
    .B(_1251_),
    .Y(_1295_));
 OA211x2_ASAP7_75t_R _4080_ (.A1(_1028_),
    .A2(_1294_),
    .B(_1295_),
    .C(_1104_),
    .Y(_1296_));
 OA21x2_ASAP7_75t_R _4081_ (.A1(_3399_),
    .A2(_1029_),
    .B(_1253_),
    .Y(_1297_));
 AO21x2_ASAP7_75t_R _4082_ (.A1(_1050_),
    .A2(_1095_),
    .B(_1297_),
    .Y(_1298_));
 OR5x2_ASAP7_75t_R _4083_ (.A(net196),
    .B(_1077_),
    .C(_1033_),
    .D(_1013_),
    .E(_1095_),
    .Y(_1299_));
 OA211x2_ASAP7_75t_R _4084_ (.A1(_1078_),
    .A2(_1298_),
    .B(_1299_),
    .C(_1094_),
    .Y(_1300_));
 AND5x2_ASAP7_75t_R _4085_ (.A(_0993_),
    .B(_1032_),
    .C(_1022_),
    .D(_1021_),
    .E(_1215_),
    .Y(_1301_));
 AO31x2_ASAP7_75t_R _4086_ (.A1(_1030_),
    .A2(_1013_),
    .A3(_1050_),
    .B(_1301_),
    .Y(_1302_));
 OA22x2_ASAP7_75t_R _4087_ (.A1(_0556_),
    .A2(_1049_),
    .B1(_1262_),
    .B2(_1122_),
    .Y(_1303_));
 XNOR2x2_ASAP7_75t_R _4088_ (.A(_1009_),
    .B(_1010_),
    .Y(_1304_));
 AND3x2_ASAP7_75t_R _4089_ (.A(_0993_),
    .B(_1032_),
    .C(_1304_),
    .Y(_1305_));
 OA31x2_ASAP7_75t_R _4090_ (.A1(_1264_),
    .A2(_1303_),
    .A3(_1305_),
    .B1(_1297_),
    .Y(_1306_));
 AND3x2_ASAP7_75t_R _4091_ (.A(_1034_),
    .B(_1013_),
    .C(_1095_),
    .Y(_1307_));
 OR5x2_ASAP7_75t_R _4092_ (.A(_1070_),
    .B(_1077_),
    .C(_1302_),
    .D(_1306_),
    .E(_1307_),
    .Y(_1308_));
 OA21x2_ASAP7_75t_R _4093_ (.A1(_1024_),
    .A2(_1304_),
    .B(net41),
    .Y(_1309_));
 OA221x2_ASAP7_75t_R _4094_ (.A1(net47),
    .A2(_1023_),
    .B1(_1309_),
    .B2(_1034_),
    .C(_1213_),
    .Y(_1310_));
 OA21x2_ASAP7_75t_R _4095_ (.A1(net41),
    .A2(_1304_),
    .B(_1115_),
    .Y(_1311_));
 OA211x2_ASAP7_75t_R _4096_ (.A1(_1024_),
    .A2(_1023_),
    .B(_1311_),
    .C(_1033_),
    .Y(_1312_));
 OR3x2_ASAP7_75t_R _4097_ (.A(_1004_),
    .B(_1310_),
    .C(_1312_),
    .Y(_1313_));
 OA211x2_ASAP7_75t_R _4098_ (.A1(_1296_),
    .A2(_1300_),
    .B(_1308_),
    .C(_1313_),
    .Y(_1314_));
 TAPCELL_ASAP7_75t_R TAP_206 ();
 INVx4_ASAP7_75t_R _4100_ (.A(_1314_),
    .Y(_3185_));
 AND2x2_ASAP7_75t_R _4101_ (.A(_0465_),
    .B(net239),
    .Y(_1315_));
 XOR2x2_ASAP7_75t_R _4102_ (.A(_1258_),
    .B(_1315_),
    .Y(_3446_));
 AO21x2_ASAP7_75t_R _4103_ (.A1(net47),
    .A2(_1223_),
    .B(_1215_),
    .Y(_1316_));
 AO21x2_ASAP7_75t_R _4104_ (.A1(_1030_),
    .A2(_1316_),
    .B(_1132_),
    .Y(_1317_));
 AO21x2_ASAP7_75t_R _4105_ (.A1(_1050_),
    .A2(_1095_),
    .B(_1070_),
    .Y(_1318_));
 AO22x2_ASAP7_75t_R _4106_ (.A1(_1070_),
    .A2(_1111_),
    .B1(_1318_),
    .B2(_1023_),
    .Y(_1319_));
 AND3x2_ASAP7_75t_R _4107_ (.A(_1104_),
    .B(_1317_),
    .C(_1319_),
    .Y(_1320_));
 OA211x2_ASAP7_75t_R _4108_ (.A1(net46),
    .A2(_1284_),
    .B(_1187_),
    .C(_1030_),
    .Y(_1321_));
 AO221x2_ASAP7_75t_R _4109_ (.A1(_1024_),
    .A2(_1075_),
    .B1(_1095_),
    .B2(_1050_),
    .C(_1132_),
    .Y(_1322_));
 OA211x2_ASAP7_75t_R _4110_ (.A1(_1098_),
    .A2(_1321_),
    .B(_1322_),
    .C(_1077_),
    .Y(_1323_));
 OA21x2_ASAP7_75t_R _4111_ (.A1(net42),
    .A2(_1033_),
    .B(_1124_),
    .Y(_1324_));
 OA211x2_ASAP7_75t_R _4112_ (.A1(_1013_),
    .A2(_1100_),
    .B(_1024_),
    .C(_1030_),
    .Y(_1325_));
 AO21x2_ASAP7_75t_R _4113_ (.A1(net46),
    .A2(_1324_),
    .B(_1325_),
    .Y(_1326_));
 AO21x2_ASAP7_75t_R _4114_ (.A1(_1030_),
    .A2(_1249_),
    .B(_1025_),
    .Y(_1327_));
 AO21x2_ASAP7_75t_R _4115_ (.A1(_1326_),
    .A2(_1327_),
    .B(_1070_),
    .Y(_1328_));
 AO21x2_ASAP7_75t_R _4116_ (.A1(_1024_),
    .A2(_1100_),
    .B(_1050_),
    .Y(_1329_));
 AO221x2_ASAP7_75t_R _4117_ (.A1(net46),
    .A2(_1075_),
    .B1(_1329_),
    .B2(_1030_),
    .C(_1098_),
    .Y(_1330_));
 OA21x2_ASAP7_75t_R _4118_ (.A1(_1025_),
    .A2(_1013_),
    .B(_1134_),
    .Y(_1331_));
 AO21x2_ASAP7_75t_R _4119_ (.A1(_1013_),
    .A2(_1075_),
    .B(_1065_),
    .Y(_1332_));
 AO221x2_ASAP7_75t_R _4120_ (.A1(_1034_),
    .A2(_1331_),
    .B1(_1332_),
    .B2(net212),
    .C(_1070_),
    .Y(_1333_));
 OA211x2_ASAP7_75t_R _4121_ (.A1(_1195_),
    .A2(_1211_),
    .B(_1333_),
    .C(_1004_),
    .Y(_1334_));
 AO221x2_ASAP7_75t_R _4122_ (.A1(_1323_),
    .A2(_1328_),
    .B1(_1330_),
    .B2(_1334_),
    .C(_0459_),
    .Y(_1335_));
 OA21x2_ASAP7_75t_R _4123_ (.A1(_1094_),
    .A2(_1320_),
    .B(_1335_),
    .Y(_1336_));
 TAPCELL_ASAP7_75t_R PHY_205 ();
 INVx4_ASAP7_75t_R _4125_ (.A(_1336_),
    .Y(_3168_));
 AND2x2_ASAP7_75t_R _4126_ (.A(_0466_),
    .B(net237),
    .Y(_1337_));
 AO21x2_ASAP7_75t_R _4127_ (.A1(_3449_),
    .A2(_1173_),
    .B(_1337_),
    .Y(_1338_));
 TAPCELL_ASAP7_75t_R PHY_204 ();
 AND3x2_ASAP7_75t_R _4129_ (.A(_3440_),
    .B(_3441_),
    .C(_1259_),
    .Y(_3476_));
 XNOR2x2_ASAP7_75t_R _4130_ (.A(_0471_),
    .B(_0704_),
    .Y(_1339_));
 AND3x2_ASAP7_75t_R _4131_ (.A(_3475_),
    .B(_3476_),
    .C(_1339_),
    .Y(_3467_));
 XNOR2x2_ASAP7_75t_R _4132_ (.A(_0470_),
    .B(_0703_),
    .Y(_1340_));
 AND3x2_ASAP7_75t_R _4133_ (.A(_3466_),
    .B(_3467_),
    .C(_1340_),
    .Y(_3460_));
 XNOR2x2_ASAP7_75t_R _4134_ (.A(_0469_),
    .B(_0702_),
    .Y(_1341_));
 AND3x2_ASAP7_75t_R _4135_ (.A(_3459_),
    .B(_3460_),
    .C(_1341_),
    .Y(_3454_));
 INVx2_ASAP7_75t_R _4136_ (.A(_0700_),
    .Y(_1342_));
 OR2x2_ASAP7_75t_R _4137_ (.A(_0459_),
    .B(_1342_),
    .Y(_1343_));
 OR2x2_ASAP7_75t_R _4138_ (.A(_1077_),
    .B(_1343_),
    .Y(_1344_));
 OR3x4_ASAP7_75t_R _4139_ (.A(_1055_),
    .B(_1132_),
    .C(_1344_),
    .Y(_3151_));
 INVx5_ASAP7_75t_R _4140_ (.A(_3151_),
    .Y(_3154_));
 AND2x2_ASAP7_75t_R _4141_ (.A(_0472_),
    .B(net227),
    .Y(_1345_));
 AND2x2_ASAP7_75t_R _4142_ (.A(_3453_),
    .B(_1173_),
    .Y(_1346_));
 NOR2x2_ASAP7_75t_R _4143_ (.A(_1345_),
    .B(_1346_),
    .Y(_3152_));
 INVx2_ASAP7_75t_R _4144_ (.A(_3152_),
    .Y(_3155_));
 OA21x2_ASAP7_75t_R _4145_ (.A1(net213),
    .A2(_1034_),
    .B(_1013_),
    .Y(_1347_));
 OA211x2_ASAP7_75t_R _4146_ (.A1(_0263_),
    .A2(_1347_),
    .B(_1239_),
    .C(_1251_),
    .Y(_1348_));
 TAPCELL_ASAP7_75t_R PHY_203 ();
 INVx3_ASAP7_75t_R _4148_ (.A(_1348_),
    .Y(_3188_));
 AND2x2_ASAP7_75t_R _4149_ (.A(_0474_),
    .B(net239),
    .Y(_1349_));
 XNOR2x2_ASAP7_75t_R _4150_ (.A(_1341_),
    .B(_1349_),
    .Y(_3457_));
 INVx2_ASAP7_75t_R _4151_ (.A(_3457_),
    .Y(_3456_));
 AND2x2_ASAP7_75t_R _4152_ (.A(_1030_),
    .B(_1239_),
    .Y(_1350_));
 AO32x2_ASAP7_75t_R _4153_ (.A1(_1033_),
    .A2(_1304_),
    .A3(_1253_),
    .B1(_1118_),
    .B2(net42),
    .Y(_1351_));
 AO21x2_ASAP7_75t_R _4154_ (.A1(net47),
    .A2(_1107_),
    .B(_1190_),
    .Y(_1352_));
 AO22x2_ASAP7_75t_R _4155_ (.A1(_1070_),
    .A2(_1351_),
    .B1(_1352_),
    .B2(_1023_),
    .Y(_1353_));
 AND2x6_ASAP7_75t_R _4156_ (.A(_1350_),
    .B(_1353_),
    .Y(_3239_));
 INVx2_ASAP7_75t_R _4157_ (.A(_3239_),
    .Y(_3156_));
 AND2x2_ASAP7_75t_R _4158_ (.A(_0475_),
    .B(net227),
    .Y(_1354_));
 AO21x2_ASAP7_75t_R _4159_ (.A1(_3459_),
    .A2(_1173_),
    .B(_1354_),
    .Y(_1355_));
 TAPCELL_ASAP7_75t_R PHY_202 ();
 OR3x2_ASAP7_75t_R _4161_ (.A(_1055_),
    .B(_1033_),
    .C(_1013_),
    .Y(_1356_));
 AND2x2_ASAP7_75t_R _4162_ (.A(_1024_),
    .B(_1124_),
    .Y(_1357_));
 OR3x2_ASAP7_75t_R _4163_ (.A(_1055_),
    .B(_1033_),
    .C(_1086_),
    .Y(_1358_));
 OA21x2_ASAP7_75t_R _4164_ (.A1(_1013_),
    .A2(_1100_),
    .B(net47),
    .Y(_1359_));
 AO221x2_ASAP7_75t_R _4165_ (.A1(_1356_),
    .A2(_1357_),
    .B1(_1358_),
    .B2(_1359_),
    .C(net196),
    .Y(_1360_));
 AO211x2_ASAP7_75t_R _4166_ (.A1(net47),
    .A2(_1086_),
    .B(_1055_),
    .C(_1070_),
    .Y(_1361_));
 AO31x2_ASAP7_75t_R _4167_ (.A1(_1024_),
    .A2(_1114_),
    .A3(_1255_),
    .B(_1361_),
    .Y(_1362_));
 AO21x2_ASAP7_75t_R _4168_ (.A1(_1360_),
    .A2(_1362_),
    .B(_1344_),
    .Y(_1363_));
 TAPCELL_ASAP7_75t_R PHY_201 ();
 AND2x2_ASAP7_75t_R _4170_ (.A(_0477_),
    .B(net237),
    .Y(_1364_));
 XOR2x2_ASAP7_75t_R _4171_ (.A(_1340_),
    .B(_1364_),
    .Y(_3463_));
 OR3x2_ASAP7_75t_R _4172_ (.A(_1033_),
    .B(_1023_),
    .C(_1027_),
    .Y(_1365_));
 AO21x2_ASAP7_75t_R _4173_ (.A1(net43),
    .A2(_1013_),
    .B(net46),
    .Y(_1366_));
 OR2x2_ASAP7_75t_R _4174_ (.A(_1070_),
    .B(_1055_),
    .Y(_1367_));
 AO21x2_ASAP7_75t_R _4175_ (.A1(_1365_),
    .A2(_1366_),
    .B(_1367_),
    .Y(_1368_));
 OA31x2_ASAP7_75t_R _4176_ (.A1(_1024_),
    .A2(_1055_),
    .A3(_1013_),
    .B1(_1124_),
    .Y(_1369_));
 OA21x2_ASAP7_75t_R _4177_ (.A1(net204),
    .A2(_1369_),
    .B(_1004_),
    .Y(_1370_));
 OR3x2_ASAP7_75t_R _4178_ (.A(net202),
    .B(_1055_),
    .C(_1013_),
    .Y(_1371_));
 AO21x2_ASAP7_75t_R _4179_ (.A1(_1025_),
    .A2(_1184_),
    .B(_1371_),
    .Y(_1372_));
 AO22x2_ASAP7_75t_R _4180_ (.A1(_1368_),
    .A2(_1370_),
    .B1(_1372_),
    .B2(_1077_),
    .Y(_1373_));
 NOR2x2_ASAP7_75t_R _4181_ (.A(_1343_),
    .B(_1373_),
    .Y(_3468_));
 INVx5_ASAP7_75t_R _4182_ (.A(_3468_),
    .Y(_3159_));
 AND2x2_ASAP7_75t_R _4183_ (.A(_0478_),
    .B(net239),
    .Y(_1374_));
 AO21x2_ASAP7_75t_R _4184_ (.A1(_3466_),
    .A2(_1173_),
    .B(_1374_),
    .Y(_1375_));
 TAPCELL_ASAP7_75t_R PHY_200 ();
 AO21x2_ASAP7_75t_R _4186_ (.A1(_1085_),
    .A2(_1270_),
    .B(_1121_),
    .Y(_1376_));
 OA211x2_ASAP7_75t_R _4187_ (.A1(_0987_),
    .A2(_1021_),
    .B(_1022_),
    .C(_1070_),
    .Y(_1377_));
 AND2x2_ASAP7_75t_R _4188_ (.A(net214),
    .B(_1377_),
    .Y(_1378_));
 AO21x2_ASAP7_75t_R _4189_ (.A1(_1083_),
    .A2(_1132_),
    .B(_1378_),
    .Y(_1379_));
 AO22x2_ASAP7_75t_R _4190_ (.A1(net212),
    .A2(_1376_),
    .B1(_1379_),
    .B2(_1025_),
    .Y(_1380_));
 AND3x2_ASAP7_75t_R _4191_ (.A(_1070_),
    .B(_1077_),
    .C(_1094_),
    .Y(_1381_));
 AND2x2_ASAP7_75t_R _4192_ (.A(_1030_),
    .B(_1381_),
    .Y(_1382_));
 AO221x2_ASAP7_75t_R _4193_ (.A1(_1034_),
    .A2(_1019_),
    .B1(_1253_),
    .B2(_1023_),
    .C(_1085_),
    .Y(_1383_));
 AND3x2_ASAP7_75t_R _4194_ (.A(net201),
    .B(_1004_),
    .C(_1094_),
    .Y(_1384_));
 AO22x2_ASAP7_75t_R _4195_ (.A1(_1034_),
    .A2(_1023_),
    .B1(_1284_),
    .B2(_1024_),
    .Y(_1385_));
 AO32x2_ASAP7_75t_R _4196_ (.A1(net212),
    .A2(net43),
    .A3(_1305_),
    .B1(_1385_),
    .B2(_1030_),
    .Y(_1386_));
 AO222x2_ASAP7_75t_R _4197_ (.A1(_1203_),
    .A2(_1381_),
    .B1(_1382_),
    .B2(_1383_),
    .C1(_1384_),
    .C2(_1386_),
    .Y(_1387_));
 AO21x2_ASAP7_75t_R _4198_ (.A1(_1350_),
    .A2(_1380_),
    .B(_1387_),
    .Y(_1388_));
 TAPCELL_ASAP7_75t_R PHY_199 ();
 INVx4_ASAP7_75t_R _4200_ (.A(_1388_),
    .Y(_3194_));
 AND2x2_ASAP7_75t_R _4201_ (.A(_0480_),
    .B(net239),
    .Y(_1389_));
 XOR2x2_ASAP7_75t_R _4202_ (.A(_1339_),
    .B(_1389_),
    .Y(_3472_));
 AO221x2_ASAP7_75t_R _4203_ (.A1(net46),
    .A2(_1075_),
    .B1(_1187_),
    .B2(_1036_),
    .C(_1077_),
    .Y(_1390_));
 AO21x2_ASAP7_75t_R _4204_ (.A1(_1023_),
    .A2(_1284_),
    .B(_1077_),
    .Y(_1391_));
 OA211x2_ASAP7_75t_R _4205_ (.A1(_1004_),
    .A2(_1184_),
    .B(_1391_),
    .C(_1030_),
    .Y(_1392_));
 OR3x2_ASAP7_75t_R _4206_ (.A(net43),
    .B(_1077_),
    .C(_1033_),
    .Y(_1393_));
 AO21x2_ASAP7_75t_R _4207_ (.A1(_1284_),
    .A2(_1393_),
    .B(net46),
    .Y(_1394_));
 AO221x2_ASAP7_75t_R _4208_ (.A1(_1013_),
    .A2(_1390_),
    .B1(_1392_),
    .B2(_1394_),
    .C(net202),
    .Y(_1395_));
 OA21x2_ASAP7_75t_R _4209_ (.A1(_1023_),
    .A2(_1213_),
    .B(_1115_),
    .Y(_1396_));
 OA22x2_ASAP7_75t_R _4210_ (.A1(net47),
    .A2(_1034_),
    .B1(_1023_),
    .B2(_1253_),
    .Y(_1397_));
 AO21x2_ASAP7_75t_R _4211_ (.A1(net43),
    .A2(_1305_),
    .B(_1070_),
    .Y(_1398_));
 AO21x2_ASAP7_75t_R _4212_ (.A1(_1030_),
    .A2(_1397_),
    .B(_1398_),
    .Y(_1399_));
 OA211x2_ASAP7_75t_R _4213_ (.A1(_1004_),
    .A2(_1396_),
    .B(_1399_),
    .C(_1094_),
    .Y(_1400_));
 AND2x6_ASAP7_75t_R _4214_ (.A(_1395_),
    .B(_1400_),
    .Y(_3244_));
 INVx3_ASAP7_75t_R _4215_ (.A(_3244_),
    .Y(_3162_));
 AND2x2_ASAP7_75t_R _4216_ (.A(_0481_),
    .B(net237),
    .Y(_1401_));
 AO21x2_ASAP7_75t_R _4217_ (.A1(_3475_),
    .A2(_1173_),
    .B(_1401_),
    .Y(_1402_));
 TAPCELL_ASAP7_75t_R PHY_198 ();
 AND2x2_ASAP7_75t_R _4219_ (.A(_1158_),
    .B(_1159_),
    .Y(_1403_));
 OA21x2_ASAP7_75t_R _4220_ (.A1(_1403_),
    .A2(_1165_),
    .B(_1160_),
    .Y(_3148_));
 AO21x2_ASAP7_75t_R _4221_ (.A1(_0418_),
    .A2(_1167_),
    .B(_0417_),
    .Y(_1404_));
 AND2x2_ASAP7_75t_R _4222_ (.A(_0416_),
    .B(_1404_),
    .Y(_3147_));
 OR2x2_ASAP7_75t_R _4223_ (.A(_1164_),
    .B(_1403_),
    .Y(_3149_));
 XOR2x2_ASAP7_75t_R _4224_ (.A(_0392_),
    .B(_0568_),
    .Y(_1405_));
 XNOR2x2_ASAP7_75t_R _4225_ (.A(net174),
    .B(_0468_),
    .Y(_1406_));
 AND3x2_ASAP7_75t_R _4226_ (.A(_3453_),
    .B(_3454_),
    .C(_1406_),
    .Y(_3494_));
 XOR2x2_ASAP7_75t_R _4227_ (.A(_0425_),
    .B(_0572_),
    .Y(_1407_));
 AND3x2_ASAP7_75t_R _4228_ (.A(_3493_),
    .B(_3494_),
    .C(_1407_),
    .Y(_3492_));
 XOR2x2_ASAP7_75t_R _4229_ (.A(_0421_),
    .B(_0571_),
    .Y(_1408_));
 AND3x2_ASAP7_75t_R _4230_ (.A(_3491_),
    .B(_3492_),
    .C(_1408_),
    .Y(_3490_));
 XOR2x2_ASAP7_75t_R _4231_ (.A(_0417_),
    .B(_0570_),
    .Y(_1409_));
 AND3x2_ASAP7_75t_R _4232_ (.A(_3489_),
    .B(_3490_),
    .C(_1409_),
    .Y(_3488_));
 XOR2x2_ASAP7_75t_R _4233_ (.A(_0410_),
    .B(_0569_),
    .Y(_1410_));
 AND3x2_ASAP7_75t_R _4234_ (.A(_3487_),
    .B(_3488_),
    .C(_1410_),
    .Y(_3486_));
 AND3x2_ASAP7_75t_R _4235_ (.A(_3485_),
    .B(_1405_),
    .C(_3486_),
    .Y(_3484_));
 XNOR2x2_ASAP7_75t_R _4236_ (.A(_0376_),
    .B(_0484_),
    .Y(_1411_));
 AND3x2_ASAP7_75t_R _4237_ (.A(_3483_),
    .B(_3484_),
    .C(_1411_),
    .Y(_3482_));
 XNOR2x2_ASAP7_75t_R _4238_ (.A(_0352_),
    .B(_0483_),
    .Y(_1412_));
 AND3x2_ASAP7_75t_R _4239_ (.A(_3481_),
    .B(_3482_),
    .C(_1412_),
    .Y(_3480_));
 OR3x2_ASAP7_75t_R _4240_ (.A(_0473_),
    .B(_0476_),
    .C(net163),
    .Y(_1413_));
 OA21x2_ASAP7_75t_R _4241_ (.A1(_0499_),
    .A2(net182),
    .B(_0498_),
    .Y(_1414_));
 OR2x2_ASAP7_75t_R _4242_ (.A(_0464_),
    .B(net179),
    .Y(_1415_));
 OA21x2_ASAP7_75t_R _4243_ (.A1(_0497_),
    .A2(net179),
    .B(_0496_),
    .Y(_1416_));
 OA21x2_ASAP7_75t_R _4244_ (.A1(_1414_),
    .A2(_1415_),
    .B(_1416_),
    .Y(_1417_));
 OR4x2_ASAP7_75t_R _4245_ (.A(_0479_),
    .B(_0482_),
    .C(net206),
    .D(net190),
    .Y(_1418_));
 OA21x2_ASAP7_75t_R _4246_ (.A1(_0495_),
    .A2(net206),
    .B(_0494_),
    .Y(_1419_));
 OR3x2_ASAP7_75t_R _4247_ (.A(_0479_),
    .B(net194),
    .C(_1419_),
    .Y(_1420_));
 OA21x2_ASAP7_75t_R _4248_ (.A1(_0493_),
    .A2(net193),
    .B(_0492_),
    .Y(_1421_));
 OA211x2_ASAP7_75t_R _4249_ (.A1(_1417_),
    .A2(_1418_),
    .B(_1420_),
    .C(_1421_),
    .Y(_1422_));
 OR4x2_ASAP7_75t_R _4250_ (.A(_0464_),
    .B(_0467_),
    .C(net181),
    .D(net176),
    .Y(_1423_));
 OR3x4_ASAP7_75t_R _4251_ (.A(_1413_),
    .B(_1418_),
    .C(_1423_),
    .Y(_1424_));
 INVx2_ASAP7_75t_R _4252_ (.A(_0701_),
    .Y(_1425_));
 OA21x2_ASAP7_75t_R _4253_ (.A1(_1425_),
    .A2(_0708_),
    .B(_0502_),
    .Y(_1426_));
 OR2x2_ASAP7_75t_R _4254_ (.A(_0458_),
    .B(_0709_),
    .Y(_1427_));
 OA21x2_ASAP7_75t_R _4255_ (.A1(_0501_),
    .A2(_0709_),
    .B(_0500_),
    .Y(_1428_));
 OA21x2_ASAP7_75t_R _4256_ (.A1(_1426_),
    .A2(_1427_),
    .B(_1428_),
    .Y(_1429_));
 OA21x2_ASAP7_75t_R _4257_ (.A1(_0491_),
    .A2(net164),
    .B(_0490_),
    .Y(_1430_));
 OA21x2_ASAP7_75t_R _4258_ (.A1(_0473_),
    .A2(_1430_),
    .B(_0489_),
    .Y(_1431_));
 OA221x2_ASAP7_75t_R _4259_ (.A1(_1413_),
    .A2(_1422_),
    .B1(_1424_),
    .B2(_1429_),
    .C(_1431_),
    .Y(_1432_));
 INVx2_ASAP7_75t_R _4260_ (.A(_0717_),
    .Y(_1433_));
 INVx2_ASAP7_75t_R _4261_ (.A(_0724_),
    .Y(_1434_));
 OR3x2_ASAP7_75t_R _4262_ (.A(_1433_),
    .B(_1434_),
    .C(_1173_),
    .Y(_1435_));
 INVx2_ASAP7_75t_R _4263_ (.A(_3479_),
    .Y(_1436_));
 INVx2_ASAP7_75t_R _4264_ (.A(_3487_),
    .Y(_1437_));
 OR3x2_ASAP7_75t_R _4265_ (.A(_1436_),
    .B(_1437_),
    .C(net195),
    .Y(_1438_));
 INVx2_ASAP7_75t_R _4266_ (.A(_0723_),
    .Y(_1439_));
 XNOR2x2_ASAP7_75t_R _4267_ (.A(_0410_),
    .B(_0569_),
    .Y(_1440_));
 OA21x2_ASAP7_75t_R _4268_ (.A1(_1439_),
    .A2(_1173_),
    .B(_1440_),
    .Y(_1441_));
 AND3x2_ASAP7_75t_R _4269_ (.A(_0723_),
    .B(net195),
    .C(_1410_),
    .Y(_1442_));
 AO211x2_ASAP7_75t_R _4270_ (.A1(_1435_),
    .A2(_1438_),
    .B(_1441_),
    .C(_1442_),
    .Y(_1443_));
 INVx2_ASAP7_75t_R _4271_ (.A(_3489_),
    .Y(_1444_));
 OR2x2_ASAP7_75t_R _4272_ (.A(_1444_),
    .B(net195),
    .Y(_1445_));
 INVx2_ASAP7_75t_R _4273_ (.A(_0485_),
    .Y(_1446_));
 INVx2_ASAP7_75t_R _4274_ (.A(_0725_),
    .Y(_1447_));
 OR3x2_ASAP7_75t_R _4275_ (.A(_1446_),
    .B(_1447_),
    .C(_1173_),
    .Y(_1448_));
 XOR2x2_ASAP7_75t_R _4276_ (.A(_0352_),
    .B(_0483_),
    .Y(_1449_));
 AO21x2_ASAP7_75t_R _4277_ (.A1(_0718_),
    .A2(net227),
    .B(_1449_),
    .Y(_1450_));
 INVx2_ASAP7_75t_R _4278_ (.A(_0718_),
    .Y(_1451_));
 OR3x2_ASAP7_75t_R _4279_ (.A(_1451_),
    .B(_1173_),
    .C(_1412_),
    .Y(_1452_));
 INVx2_ASAP7_75t_R _4280_ (.A(_0719_),
    .Y(_1453_));
 OR2x2_ASAP7_75t_R _4281_ (.A(_1453_),
    .B(_1173_),
    .Y(_1454_));
 INVx2_ASAP7_75t_R _4282_ (.A(_3481_),
    .Y(_1455_));
 OR2x2_ASAP7_75t_R _4283_ (.A(_1455_),
    .B(net227),
    .Y(_1456_));
 AO222x2_ASAP7_75t_R _4284_ (.A1(_1445_),
    .A2(_1448_),
    .B1(_1450_),
    .B2(_1452_),
    .C1(_1454_),
    .C2(_1456_),
    .Y(_1457_));
 OR3x4_ASAP7_75t_R _4285_ (.A(_1432_),
    .B(_1443_),
    .C(_1457_),
    .Y(_1458_));
 INVx2_ASAP7_75t_R _4286_ (.A(_0727_),
    .Y(_1459_));
 OR2x2_ASAP7_75t_R _4287_ (.A(_1459_),
    .B(_1173_),
    .Y(_1460_));
 INVx2_ASAP7_75t_R _4288_ (.A(_3491_),
    .Y(_1461_));
 OR2x2_ASAP7_75t_R _4289_ (.A(_1461_),
    .B(net195),
    .Y(_1462_));
 INVx2_ASAP7_75t_R _4290_ (.A(_0726_),
    .Y(_1463_));
 XNOR2x2_ASAP7_75t_R _4291_ (.A(_0421_),
    .B(_0571_),
    .Y(_1464_));
 OA21x2_ASAP7_75t_R _4292_ (.A1(_1463_),
    .A2(_1173_),
    .B(_1464_),
    .Y(_1465_));
 AND3x2_ASAP7_75t_R _4293_ (.A(_0726_),
    .B(net195),
    .C(_1408_),
    .Y(_1466_));
 AO211x2_ASAP7_75t_R _4294_ (.A1(_1460_),
    .A2(_1462_),
    .B(_1465_),
    .C(_1466_),
    .Y(_1467_));
 AND3x2_ASAP7_75t_R _4295_ (.A(_3493_),
    .B(_1173_),
    .C(_1407_),
    .Y(_1468_));
 XNOR2x2_ASAP7_75t_R _4296_ (.A(_0425_),
    .B(_0572_),
    .Y(_1469_));
 XNOR2x2_ASAP7_75t_R _4297_ (.A(_0488_),
    .B(_1469_),
    .Y(_1470_));
 AND3x2_ASAP7_75t_R _4298_ (.A(_0728_),
    .B(net195),
    .C(_1470_),
    .Y(_1471_));
 NOR2x2_ASAP7_75t_R _4299_ (.A(_1468_),
    .B(_1471_),
    .Y(_1472_));
 INVx2_ASAP7_75t_R _4300_ (.A(_3485_),
    .Y(_1473_));
 INVx2_ASAP7_75t_R _4301_ (.A(_1405_),
    .Y(_1474_));
 OR3x2_ASAP7_75t_R _4302_ (.A(_1473_),
    .B(net227),
    .C(_1474_),
    .Y(_1475_));
 INVx2_ASAP7_75t_R _4303_ (.A(_0721_),
    .Y(_1476_));
 XNOR2x2_ASAP7_75t_R _4304_ (.A(_1476_),
    .B(_1405_),
    .Y(_1477_));
 NAND3x2_ASAP7_75t_R _4305_ (.B(net195),
    .C(_1477_),
    .Y(_1478_),
    .A(_0722_));
 XOR2x2_ASAP7_75t_R _4306_ (.A(_0376_),
    .B(_0484_),
    .Y(_1479_));
 AO21x2_ASAP7_75t_R _4307_ (.A1(_0486_),
    .A2(net227),
    .B(_1479_),
    .Y(_1480_));
 INVx2_ASAP7_75t_R _4308_ (.A(_0486_),
    .Y(_1481_));
 OR3x2_ASAP7_75t_R _4309_ (.A(_1481_),
    .B(_1173_),
    .C(_1411_),
    .Y(_1482_));
 INVx2_ASAP7_75t_R _4310_ (.A(_3483_),
    .Y(_1483_));
 OR3x2_ASAP7_75t_R _4311_ (.A(_1171_),
    .B(_1483_),
    .C(_1172_),
    .Y(_1484_));
 INVx2_ASAP7_75t_R _4312_ (.A(_0720_),
    .Y(_1485_));
 OR3x2_ASAP7_75t_R _4313_ (.A(_0567_),
    .B(_1485_),
    .C(_1172_),
    .Y(_1486_));
 XOR2x2_ASAP7_75t_R _4314_ (.A(_0453_),
    .B(_3145_),
    .Y(_1487_));
 OR3x2_ASAP7_75t_R _4315_ (.A(_0567_),
    .B(_1483_),
    .C(_1487_),
    .Y(_1488_));
 OR3x2_ASAP7_75t_R _4316_ (.A(_1171_),
    .B(_1485_),
    .C(_1487_),
    .Y(_1489_));
 AND4x2_ASAP7_75t_R _4317_ (.A(_1484_),
    .B(_1486_),
    .C(_1488_),
    .D(_1489_),
    .Y(_1490_));
 AO221x2_ASAP7_75t_R _4318_ (.A1(_1475_),
    .A2(_1478_),
    .B1(_1480_),
    .B2(_1482_),
    .C(_1490_),
    .Y(_1491_));
 INVx2_ASAP7_75t_R _4319_ (.A(_0712_),
    .Y(_1492_));
 OA21x2_ASAP7_75t_R _4320_ (.A1(_1492_),
    .A2(_1173_),
    .B(_1406_),
    .Y(_1493_));
 TAPCELL_ASAP7_75t_R PHY_197 ();
 XOR2x2_ASAP7_75t_R _4322_ (.A(net175),
    .B(_0468_),
    .Y(_1495_));
 AND3x4_ASAP7_75t_R _4323_ (.A(_0712_),
    .B(net195),
    .C(_1495_),
    .Y(_1496_));
 NOR2x2_ASAP7_75t_R _4324_ (.A(_1493_),
    .B(_1496_),
    .Y(_1497_));
 OR3x4_ASAP7_75t_R _4325_ (.A(_0285_),
    .B(_0708_),
    .C(_1427_),
    .Y(_1498_));
 NOR2x2_ASAP7_75t_R _4326_ (.A(_1424_),
    .B(_1498_),
    .Y(_1499_));
 INVx2_ASAP7_75t_R _4327_ (.A(_0487_),
    .Y(_1500_));
 XNOR2x2_ASAP7_75t_R _4328_ (.A(_0417_),
    .B(_0570_),
    .Y(_1501_));
 OA21x2_ASAP7_75t_R _4329_ (.A1(_1500_),
    .A2(_1173_),
    .B(_1501_),
    .Y(_1502_));
 AND3x2_ASAP7_75t_R _4330_ (.A(_0487_),
    .B(net227),
    .C(_1409_),
    .Y(_1503_));
 OR3x2_ASAP7_75t_R _4331_ (.A(_1499_),
    .B(_1502_),
    .C(_1503_),
    .Y(_1504_));
 OR5x2_ASAP7_75t_R _4332_ (.A(_1467_),
    .B(_1472_),
    .C(_1491_),
    .D(_1497_),
    .E(_1504_),
    .Y(_1505_));
 OR2x4_ASAP7_75t_R _4333_ (.A(_0485_),
    .B(_1173_),
    .Y(_1506_));
 OA21x2_ASAP7_75t_R _4334_ (.A1(_1458_),
    .A2(_1505_),
    .B(_1506_),
    .Y(_1507_));
 CKINVDCx20_ASAP7_75t_R _4335_ (.A(net38),
    .Y(_1508_));
 TAPCELL_ASAP7_75t_R PHY_196 ();
 TAPCELL_ASAP7_75t_R PHY_195 ();
 TAPCELL_ASAP7_75t_R PHY_194 ();
 TAPCELL_ASAP7_75t_R PHY_193 ();
 TAPCELL_ASAP7_75t_R PHY_192 ();
 TAPCELL_ASAP7_75t_R PHY_191 ();
 TAPCELL_ASAP7_75t_R PHY_190 ();
 OA21x2_ASAP7_75t_R _4343_ (.A1(_0009_),
    .A2(net184),
    .B(_0008_),
    .Y(_1515_));
 OA21x2_ASAP7_75t_R _4344_ (.A1(_0464_),
    .A2(_1515_),
    .B(_0007_),
    .Y(_1516_));
 OA21x2_ASAP7_75t_R _4345_ (.A1(_0458_),
    .A2(_0012_),
    .B(_0011_),
    .Y(_1517_));
 OA21x2_ASAP7_75t_R _4346_ (.A1(_0709_),
    .A2(_1517_),
    .B(_0010_),
    .Y(_1518_));
 OA21x2_ASAP7_75t_R _4347_ (.A1(_1423_),
    .A2(_1518_),
    .B(_0006_),
    .Y(_1519_));
 OA21x2_ASAP7_75t_R _4348_ (.A1(net177),
    .A2(_1516_),
    .B(_1519_),
    .Y(_1520_));
 OA21x2_ASAP7_75t_R _4349_ (.A1(_0482_),
    .A2(_1520_),
    .B(_0005_),
    .Y(_1521_));
 OA21x2_ASAP7_75t_R _4350_ (.A1(net208),
    .A2(_1521_),
    .B(_0004_),
    .Y(_1522_));
 OA21x2_ASAP7_75t_R _4351_ (.A1(_0479_),
    .A2(_1522_),
    .B(_0003_),
    .Y(_1523_));
 OA21x2_ASAP7_75t_R _4352_ (.A1(net191),
    .A2(_1523_),
    .B(_0002_),
    .Y(_1524_));
 OA21x2_ASAP7_75t_R _4353_ (.A1(_0001_),
    .A2(net166),
    .B(_0000_),
    .Y(_1525_));
 OR2x2_ASAP7_75t_R _4354_ (.A(_1493_),
    .B(_1496_),
    .Y(_1526_));
 OA211x2_ASAP7_75t_R _4355_ (.A1(_0473_),
    .A2(_1525_),
    .B(_1526_),
    .C(_0713_),
    .Y(_1527_));
 OA21x2_ASAP7_75t_R _4356_ (.A1(_1413_),
    .A2(_1524_),
    .B(_1527_),
    .Y(_3510_));
 AO21x2_ASAP7_75t_R _4357_ (.A1(_0723_),
    .A2(net195),
    .B(_1410_),
    .Y(_1528_));
 OR3x2_ASAP7_75t_R _4358_ (.A(_1439_),
    .B(net209),
    .C(_1440_),
    .Y(_1529_));
 AND2x2_ASAP7_75t_R _4359_ (.A(_1528_),
    .B(_1529_),
    .Y(_1530_));
 AND2x2_ASAP7_75t_R _4360_ (.A(_0724_),
    .B(net195),
    .Y(_1531_));
 AO21x2_ASAP7_75t_R _4361_ (.A1(_3487_),
    .A2(net209),
    .B(_1531_),
    .Y(_1532_));
 TAPCELL_ASAP7_75t_R PHY_189 ();
 TAPCELL_ASAP7_75t_R PHY_188 ();
 AO21x2_ASAP7_75t_R _4364_ (.A1(_0487_),
    .A2(net195),
    .B(_1409_),
    .Y(_1534_));
 OR3x4_ASAP7_75t_R _4365_ (.A(_1500_),
    .B(net209),
    .C(_1501_),
    .Y(_1535_));
 AND2x2_ASAP7_75t_R _4366_ (.A(_3489_),
    .B(net209),
    .Y(_1536_));
 AO21x2_ASAP7_75t_R _4367_ (.A1(_0725_),
    .A2(net195),
    .B(_1536_),
    .Y(_3505_));
 AND3x2_ASAP7_75t_R _4368_ (.A(_1534_),
    .B(_1535_),
    .C(_3505_),
    .Y(_1537_));
 AND2x2_ASAP7_75t_R _4369_ (.A(_0727_),
    .B(net195),
    .Y(_1538_));
 AND2x2_ASAP7_75t_R _4370_ (.A(_3491_),
    .B(net209),
    .Y(_1539_));
 AO21x2_ASAP7_75t_R _4371_ (.A1(_0726_),
    .A2(net195),
    .B(_1408_),
    .Y(_1540_));
 OR3x2_ASAP7_75t_R _4372_ (.A(_1463_),
    .B(net209),
    .C(_1464_),
    .Y(_1541_));
 OA211x2_ASAP7_75t_R _4373_ (.A1(_1538_),
    .A2(_1539_),
    .B(_1540_),
    .C(_1541_),
    .Y(_1542_));
 TAPCELL_ASAP7_75t_R PHY_187 ();
 OR2x2_ASAP7_75t_R _4375_ (.A(_1468_),
    .B(_1471_),
    .Y(_1544_));
 AND2x2_ASAP7_75t_R _4376_ (.A(_1544_),
    .B(_3510_),
    .Y(_3508_));
 AND2x2_ASAP7_75t_R _4377_ (.A(_1542_),
    .B(_3508_),
    .Y(_3506_));
 AND2x2_ASAP7_75t_R _4378_ (.A(_1537_),
    .B(_3506_),
    .Y(_3504_));
 AND3x2_ASAP7_75t_R _4379_ (.A(_1530_),
    .B(_1532_),
    .C(_3504_),
    .Y(_3502_));
 AND3x2_ASAP7_75t_R _4380_ (.A(_3485_),
    .B(net209),
    .C(_1405_),
    .Y(_1545_));
 AND3x2_ASAP7_75t_R _4381_ (.A(_0722_),
    .B(net195),
    .C(_1477_),
    .Y(_1546_));
 OA21x2_ASAP7_75t_R _4382_ (.A1(_1481_),
    .A2(net209),
    .B(_1411_),
    .Y(_1547_));
 AND3x2_ASAP7_75t_R _4383_ (.A(_0486_),
    .B(net162),
    .C(_1479_),
    .Y(_1548_));
 INVx2_ASAP7_75t_R _4384_ (.A(_1490_),
    .Y(_3499_));
 OA221x2_ASAP7_75t_R _4385_ (.A1(_1545_),
    .A2(_1546_),
    .B1(_1547_),
    .B2(_1548_),
    .C(_3499_),
    .Y(_1549_));
 AND2x2_ASAP7_75t_R _4386_ (.A(_1549_),
    .B(_3502_),
    .Y(_3498_));
 OA21x2_ASAP7_75t_R _4387_ (.A1(_1451_),
    .A2(net209),
    .B(_1412_),
    .Y(_1550_));
 AND3x2_ASAP7_75t_R _4388_ (.A(_0718_),
    .B(net162),
    .C(_1449_),
    .Y(_1551_));
 OR2x2_ASAP7_75t_R _4389_ (.A(_1550_),
    .B(_1551_),
    .Y(_1552_));
 NAND2x2_ASAP7_75t_R _4390_ (.A(_1454_),
    .B(_1456_),
    .Y(_3497_));
 AND3x2_ASAP7_75t_R _4391_ (.A(_1552_),
    .B(_3497_),
    .C(_3498_),
    .Y(_3496_));
 OR2x2_ASAP7_75t_R _4392_ (.A(_1545_),
    .B(_1546_),
    .Y(_1553_));
 AND2x2_ASAP7_75t_R _4393_ (.A(_1553_),
    .B(_3502_),
    .Y(_3500_));
 TAPCELL_ASAP7_75t_R PHY_186 ();
 TAPCELL_ASAP7_75t_R PHY_185 ();
 TAPCELL_ASAP7_75t_R PHY_184 ();
 TAPCELL_ASAP7_75t_R PHY_183 ();
 TAPCELL_ASAP7_75t_R PHY_182 ();
 TAPCELL_ASAP7_75t_R PHY_181 ();
 TAPCELL_ASAP7_75t_R PHY_180 ();
 XOR2x2_ASAP7_75t_R _4401_ (.A(_0023_),
    .B(net167),
    .Y(_1560_));
 AND2x2_ASAP7_75t_R _4402_ (.A(_3457_),
    .B(_1508_),
    .Y(_1561_));
 AO21x2_ASAP7_75t_R _4403_ (.A1(net39),
    .A2(_1560_),
    .B(_1561_),
    .Y(_3511_));
 INVx2_ASAP7_75t_R _4404_ (.A(_3511_),
    .Y(_3512_));
 TAPCELL_ASAP7_75t_R PHY_179 ();
 OR2x2_ASAP7_75t_R _4406_ (.A(_1355_),
    .B(net39),
    .Y(_1563_));
 OA21x2_ASAP7_75t_R _4407_ (.A1(_0026_),
    .A2(_1508_),
    .B(_1563_),
    .Y(_1564_));
 TAPCELL_ASAP7_75t_R PHY_178 ();
 TAPCELL_ASAP7_75t_R PHY_177 ();
 XNOR2x2_ASAP7_75t_R _4410_ (.A(_0028_),
    .B(net192),
    .Y(_1566_));
 OR2x2_ASAP7_75t_R _4411_ (.A(_1508_),
    .B(_1566_),
    .Y(_1567_));
 OA21x2_ASAP7_75t_R _4412_ (.A1(_3463_),
    .A2(net39),
    .B(_1567_),
    .Y(_1568_));
 TAPCELL_ASAP7_75t_R PHY_176 ();
 OR2x2_ASAP7_75t_R _4414_ (.A(_1375_),
    .B(net39),
    .Y(_1569_));
 OA21x2_ASAP7_75t_R _4415_ (.A1(_0030_),
    .A2(_1508_),
    .B(_1569_),
    .Y(_1570_));
 TAPCELL_ASAP7_75t_R PHY_175 ();
 XNOR2x2_ASAP7_75t_R _4417_ (.A(_0033_),
    .B(net207),
    .Y(_1571_));
 OR2x2_ASAP7_75t_R _4418_ (.A(_1508_),
    .B(_1571_),
    .Y(_1572_));
 OA21x2_ASAP7_75t_R _4419_ (.A1(_3472_),
    .A2(net39),
    .B(_1572_),
    .Y(_1573_));
 TAPCELL_ASAP7_75t_R PHY_174 ();
 OR2x2_ASAP7_75t_R _4421_ (.A(_1402_),
    .B(net39),
    .Y(_1574_));
 OA21x2_ASAP7_75t_R _4422_ (.A1(_0035_),
    .A2(_1508_),
    .B(_1574_),
    .Y(_1575_));
 TAPCELL_ASAP7_75t_R PHY_173 ();
 XNOR2x2_ASAP7_75t_R _4424_ (.A(_0038_),
    .B(net178),
    .Y(_1576_));
 OR2x2_ASAP7_75t_R _4425_ (.A(_1508_),
    .B(_1576_),
    .Y(_1577_));
 OA21x2_ASAP7_75t_R _4426_ (.A1(_3437_),
    .A2(net39),
    .B(_1577_),
    .Y(_1578_));
 TAPCELL_ASAP7_75t_R PHY_172 ();
 OR2x2_ASAP7_75t_R _4428_ (.A(_1293_),
    .B(net39),
    .Y(_1579_));
 OA21x2_ASAP7_75t_R _4429_ (.A1(_0040_),
    .A2(_1508_),
    .B(_1579_),
    .Y(_1580_));
 TAPCELL_ASAP7_75t_R PHY_171 ();
 XNOR2x2_ASAP7_75t_R _4431_ (.A(_0043_),
    .B(net183),
    .Y(_1581_));
 AND2x2_ASAP7_75t_R _4432_ (.A(net39),
    .B(_1581_),
    .Y(_1582_));
 AO21x2_ASAP7_75t_R _4433_ (.A1(_3446_),
    .A2(_1508_),
    .B(_1582_),
    .Y(_1583_));
 TAPCELL_ASAP7_75t_R PHY_170 ();
 OR2x2_ASAP7_75t_R _4435_ (.A(_1338_),
    .B(net39),
    .Y(_1584_));
 OA21x2_ASAP7_75t_R _4436_ (.A1(_0045_),
    .A2(_1508_),
    .B(_1584_),
    .Y(_1585_));
 TAPCELL_ASAP7_75t_R PHY_169 ();
 XNOR2x2_ASAP7_75t_R _4438_ (.A(_0048_),
    .B(_0709_),
    .Y(_1586_));
 OR2x2_ASAP7_75t_R _4439_ (.A(_1508_),
    .B(_1586_),
    .Y(_1587_));
 OA21x2_ASAP7_75t_R _4440_ (.A1(_3430_),
    .A2(net39),
    .B(_1587_),
    .Y(_1588_));
 TAPCELL_ASAP7_75t_R PHY_168 ();
 OR2x2_ASAP7_75t_R _4442_ (.A(_1238_),
    .B(net39),
    .Y(_1589_));
 OA21x2_ASAP7_75t_R _4443_ (.A1(_0050_),
    .A2(_1508_),
    .B(_1589_),
    .Y(_1590_));
 TAPCELL_ASAP7_75t_R PHY_167 ();
 OR2x2_ASAP7_75t_R _4445_ (.A(_1183_),
    .B(net39),
    .Y(_1591_));
 OA21x2_ASAP7_75t_R _4446_ (.A1(_0053_),
    .A2(_1508_),
    .B(_1591_),
    .Y(_1592_));
 TAPCELL_ASAP7_75t_R PHY_166 ();
 INVx2_ASAP7_75t_R _4448_ (.A(_3408_),
    .Y(_3406_));
 AND2x2_ASAP7_75t_R _4449_ (.A(_0285_),
    .B(net39),
    .Y(_1593_));
 AO21x2_ASAP7_75t_R _4450_ (.A1(_3408_),
    .A2(_1508_),
    .B(_1593_),
    .Y(_1594_));
 TAPCELL_ASAP7_75t_R PHY_165 ();
 INVx2_ASAP7_75t_R _4452_ (.A(_1594_),
    .Y(_3542_));
 INVx2_ASAP7_75t_R _4453_ (.A(_0733_),
    .Y(_1595_));
 OR2x2_ASAP7_75t_R _4454_ (.A(_1458_),
    .B(_1505_),
    .Y(_1596_));
 AND2x4_ASAP7_75t_R _4455_ (.A(_1446_),
    .B(net162),
    .Y(_1597_));
 AO21x2_ASAP7_75t_R _4456_ (.A1(_1595_),
    .A2(_1596_),
    .B(_1597_),
    .Y(_1598_));
 TAPCELL_ASAP7_75t_R PHY_164 ();
 AND2x2_ASAP7_75t_R _4458_ (.A(_1450_),
    .B(_1452_),
    .Y(_1600_));
 OR4x2_ASAP7_75t_R _4459_ (.A(_0485_),
    .B(_1453_),
    .C(net209),
    .D(_1600_),
    .Y(_1601_));
 INVx2_ASAP7_75t_R _4460_ (.A(_0734_),
    .Y(_1602_));
 AO21x2_ASAP7_75t_R _4461_ (.A1(_1450_),
    .A2(_1452_),
    .B(_1602_),
    .Y(_1603_));
 OR3x2_ASAP7_75t_R _4462_ (.A(_0734_),
    .B(_1550_),
    .C(_1551_),
    .Y(_1604_));
 AO221x2_ASAP7_75t_R _4463_ (.A1(_1446_),
    .A2(net162),
    .B1(_1603_),
    .B2(_1604_),
    .C(_0014_),
    .Y(_1605_));
 NAND2x2_ASAP7_75t_R _4464_ (.A(_1601_),
    .B(_1605_),
    .Y(_1606_));
 INVx2_ASAP7_75t_R _4465_ (.A(_0022_),
    .Y(_1607_));
 TAPCELL_ASAP7_75t_R PHY_163 ();
 NOR3x2_ASAP7_75t_R _4467_ (.B(_1493_),
    .C(_1496_),
    .Y(_1609_),
    .A(_0021_));
 OA21x2_ASAP7_75t_R _4468_ (.A1(_1493_),
    .A2(_1496_),
    .B(_0021_),
    .Y(_1610_));
 NOR2x2_ASAP7_75t_R _4469_ (.A(_1609_),
    .B(_1610_),
    .Y(_1611_));
 AND2x2_ASAP7_75t_R _4470_ (.A(_1607_),
    .B(_1611_),
    .Y(_1612_));
 AND3x2_ASAP7_75t_R _4471_ (.A(net39),
    .B(_1606_),
    .C(_1612_),
    .Y(_1613_));
 AND2x2_ASAP7_75t_R _4472_ (.A(_3155_),
    .B(_1526_),
    .Y(_1614_));
 INVx2_ASAP7_75t_R _4473_ (.A(_1614_),
    .Y(_1615_));
 OA21x2_ASAP7_75t_R _4474_ (.A1(_1458_),
    .A2(_1505_),
    .B(_1601_),
    .Y(_1616_));
 NOR2x2_ASAP7_75t_R _4475_ (.A(_1615_),
    .B(_1616_),
    .Y(_1617_));
 NOR2x2_ASAP7_75t_R _4476_ (.A(_1443_),
    .B(net39),
    .Y(_1618_));
 INVx2_ASAP7_75t_R _4477_ (.A(_0737_),
    .Y(_1619_));
 XNOR2x2_ASAP7_75t_R _4478_ (.A(_1619_),
    .B(_1530_),
    .Y(_1620_));
 OR3x4_ASAP7_75t_R _4479_ (.A(_0013_),
    .B(_0017_),
    .C(_1620_),
    .Y(_1621_));
 NOR2x2_ASAP7_75t_R _4480_ (.A(_1508_),
    .B(_1621_),
    .Y(_1622_));
 OR4x2_ASAP7_75t_R _4481_ (.A(_0042_),
    .B(_0047_),
    .C(_0745_),
    .D(_0744_),
    .Y(_1623_));
 INVx2_ASAP7_75t_R _4482_ (.A(_0749_),
    .Y(_1624_));
 OA21x2_ASAP7_75t_R _4483_ (.A1(_1624_),
    .A2(_0747_),
    .B(_0054_),
    .Y(_1625_));
 OA21x2_ASAP7_75t_R _4484_ (.A1(_0052_),
    .A2(_1625_),
    .B(_0051_),
    .Y(_1626_));
 OA21x2_ASAP7_75t_R _4485_ (.A1(_0746_),
    .A2(_1626_),
    .B(_0049_),
    .Y(_1627_));
 OA21x2_ASAP7_75t_R _4486_ (.A1(_0046_),
    .A2(_0745_),
    .B(_0044_),
    .Y(_1628_));
 OA21x2_ASAP7_75t_R _4487_ (.A1(_0042_),
    .A2(_1628_),
    .B(_0041_),
    .Y(_1629_));
 OA21x2_ASAP7_75t_R _4488_ (.A1(_0036_),
    .A2(_0743_),
    .B(_0034_),
    .Y(_1630_));
 OA21x2_ASAP7_75t_R _4489_ (.A1(_0032_),
    .A2(_1630_),
    .B(_0031_),
    .Y(_1631_));
 OA211x2_ASAP7_75t_R _4490_ (.A1(net169),
    .A2(_0741_),
    .B(_0029_),
    .C(_0024_),
    .Y(_1632_));
 OA21x2_ASAP7_75t_R _4491_ (.A1(_0742_),
    .A2(_1631_),
    .B(_1632_),
    .Y(_1633_));
 OA211x2_ASAP7_75t_R _4492_ (.A1(_0744_),
    .A2(_1629_),
    .B(_1633_),
    .C(_0039_),
    .Y(_1634_));
 OA21x2_ASAP7_75t_R _4493_ (.A1(_1623_),
    .A2(_1627_),
    .B(_1634_),
    .Y(_1635_));
 AO21x2_ASAP7_75t_R _4494_ (.A1(_0027_),
    .A2(_0741_),
    .B(net172),
    .Y(_1636_));
 OR4x2_ASAP7_75t_R _4495_ (.A(_0032_),
    .B(_0037_),
    .C(net187),
    .D(_0742_),
    .Y(_1637_));
 OR4x2_ASAP7_75t_R _4496_ (.A(net169),
    .B(_0027_),
    .C(_0052_),
    .D(_0748_),
    .Y(_1638_));
 OR4x2_ASAP7_75t_R _4497_ (.A(_0747_),
    .B(_0746_),
    .C(_1623_),
    .D(_1638_),
    .Y(_1639_));
 NOR2x2_ASAP7_75t_R _4498_ (.A(_1637_),
    .B(_1639_),
    .Y(_1640_));
 AO221x2_ASAP7_75t_R _4499_ (.A1(_0024_),
    .A2(_1636_),
    .B1(_1637_),
    .B2(_1633_),
    .C(_1640_),
    .Y(_1641_));
 NOR2x2_ASAP7_75t_R _4500_ (.A(_1635_),
    .B(_1641_),
    .Y(_1642_));
 AND4x2_ASAP7_75t_R _4501_ (.A(_1542_),
    .B(_1544_),
    .C(_1549_),
    .D(_1537_),
    .Y(_1643_));
 AND3x2_ASAP7_75t_R _4502_ (.A(_1508_),
    .B(_1642_),
    .C(_1643_),
    .Y(_1644_));
 TAPCELL_ASAP7_75t_R PHY_162 ();
 INVx2_ASAP7_75t_R _4504_ (.A(_0488_),
    .Y(_1646_));
 OA21x2_ASAP7_75t_R _4505_ (.A1(_1646_),
    .A2(net209),
    .B(_1469_),
    .Y(_1647_));
 AND3x2_ASAP7_75t_R _4506_ (.A(_0488_),
    .B(net162),
    .C(_1407_),
    .Y(_1648_));
 NOR3x2_ASAP7_75t_R _4507_ (.B(_1647_),
    .C(_1648_),
    .Y(_1649_),
    .A(_0740_));
 OA21x2_ASAP7_75t_R _4508_ (.A1(_1647_),
    .A2(_1648_),
    .B(_0740_),
    .Y(_1650_));
 NOR3x2_ASAP7_75t_R _4509_ (.B(_1649_),
    .C(_1650_),
    .Y(_1651_),
    .A(_0020_));
 INVx2_ASAP7_75t_R _4510_ (.A(_0019_),
    .Y(_1652_));
 INVx2_ASAP7_75t_R _4511_ (.A(_0018_),
    .Y(_1653_));
 OR3x2_ASAP7_75t_R _4512_ (.A(_0738_),
    .B(_1502_),
    .C(_1503_),
    .Y(_1654_));
 INVx2_ASAP7_75t_R _4513_ (.A(_0738_),
    .Y(_1655_));
 AO21x2_ASAP7_75t_R _4514_ (.A1(_1534_),
    .A2(_1535_),
    .B(_1655_),
    .Y(_1656_));
 AND3x2_ASAP7_75t_R _4515_ (.A(_1653_),
    .B(_1654_),
    .C(_1656_),
    .Y(_1657_));
 OA21x2_ASAP7_75t_R _4516_ (.A1(_1547_),
    .A2(_1548_),
    .B(_0735_),
    .Y(_1658_));
 INVx2_ASAP7_75t_R _4517_ (.A(_0735_),
    .Y(_1659_));
 AND3x2_ASAP7_75t_R _4518_ (.A(_1659_),
    .B(_1480_),
    .C(_1482_),
    .Y(_1660_));
 XNOR2x2_ASAP7_75t_R _4519_ (.A(_0736_),
    .B(_1405_),
    .Y(_1661_));
 OA21x2_ASAP7_75t_R _4520_ (.A1(_1476_),
    .A2(net209),
    .B(_1661_),
    .Y(_1662_));
 INVx2_ASAP7_75t_R _4521_ (.A(_0736_),
    .Y(_1663_));
 XNOR2x2_ASAP7_75t_R _4522_ (.A(_1663_),
    .B(_1405_),
    .Y(_1664_));
 AND3x2_ASAP7_75t_R _4523_ (.A(_0721_),
    .B(net162),
    .C(_1664_),
    .Y(_1665_));
 INVx2_ASAP7_75t_R _4524_ (.A(_0015_),
    .Y(_1666_));
 INVx2_ASAP7_75t_R _4525_ (.A(_0016_),
    .Y(_1667_));
 OA211x2_ASAP7_75t_R _4526_ (.A1(_1662_),
    .A2(_1665_),
    .B(_1666_),
    .C(_1667_),
    .Y(_1668_));
 OA21x2_ASAP7_75t_R _4527_ (.A1(_1658_),
    .A2(_1660_),
    .B(_1668_),
    .Y(_1669_));
 OR2x4_ASAP7_75t_R _4528_ (.A(_1465_),
    .B(_1466_),
    .Y(_1670_));
 XOR2x2_ASAP7_75t_R _4529_ (.A(_0739_),
    .B(_1670_),
    .Y(_1671_));
 AND4x2_ASAP7_75t_R _4530_ (.A(_1652_),
    .B(_1657_),
    .C(_1669_),
    .D(_1671_),
    .Y(_1672_));
 AND4x2_ASAP7_75t_R _4531_ (.A(net39),
    .B(_1642_),
    .C(_1651_),
    .D(_1672_),
    .Y(_1673_));
 OA222x2_ASAP7_75t_R _4532_ (.A1(_1613_),
    .A2(_1617_),
    .B1(_1618_),
    .B2(_1622_),
    .C1(_1644_),
    .C2(_1673_),
    .Y(_1674_));
 TAPCELL_ASAP7_75t_R PHY_161 ();
 OR2x6_ASAP7_75t_R _4534_ (.A(_1598_),
    .B(_1674_),
    .Y(_1676_));
 CKINVDCx20_ASAP7_75t_R _4535_ (.A(_1676_),
    .Y(_1677_));
 TAPCELL_ASAP7_75t_R PHY_160 ();
 TAPCELL_ASAP7_75t_R PHY_159 ();
 TAPCELL_ASAP7_75t_R PHY_158 ();
 TAPCELL_ASAP7_75t_R PHY_157 ();
 TAPCELL_ASAP7_75t_R PHY_156 ();
 TAPCELL_ASAP7_75t_R PHY_155 ();
 TAPCELL_ASAP7_75t_R PHY_154 ();
 TAPCELL_ASAP7_75t_R PHY_153 ();
 TAPCELL_ASAP7_75t_R PHY_152 ();
 AND2x2_ASAP7_75t_R _4545_ (.A(_1592_),
    .B(net225),
    .Y(_1686_));
 AO21x2_ASAP7_75t_R _4546_ (.A1(_0056_),
    .A2(_1677_),
    .B(_1686_),
    .Y(_3546_));
 XNOR2x2_ASAP7_75t_R _4547_ (.A(_0060_),
    .B(_0746_),
    .Y(_1687_));
 OR2x2_ASAP7_75t_R _4548_ (.A(_1588_),
    .B(_1677_),
    .Y(_1688_));
 OA21x2_ASAP7_75t_R _4549_ (.A1(net221),
    .A2(_1687_),
    .B(_1688_),
    .Y(_3547_));
 AND2x2_ASAP7_75t_R _4550_ (.A(_1590_),
    .B(net225),
    .Y(_1689_));
 AO21x2_ASAP7_75t_R _4551_ (.A1(_0061_),
    .A2(_1677_),
    .B(_1689_),
    .Y(_3548_));
 XNOR2x2_ASAP7_75t_R _4552_ (.A(_0067_),
    .B(net220),
    .Y(_1690_));
 OR2x2_ASAP7_75t_R _4553_ (.A(_1578_),
    .B(_1677_),
    .Y(_1691_));
 OA21x2_ASAP7_75t_R _4554_ (.A1(net225),
    .A2(_1690_),
    .B(_1691_),
    .Y(_3549_));
 INVx2_ASAP7_75t_R _4555_ (.A(_1580_),
    .Y(_3183_));
 XNOR2x2_ASAP7_75t_R _4556_ (.A(_0070_),
    .B(net232),
    .Y(_1692_));
 OR2x2_ASAP7_75t_R _4557_ (.A(_1583_),
    .B(_1677_),
    .Y(_1693_));
 OA21x2_ASAP7_75t_R _4558_ (.A1(net225),
    .A2(_1692_),
    .B(_1693_),
    .Y(_3551_));
 INVx2_ASAP7_75t_R _4559_ (.A(_1585_),
    .Y(_3186_));
 OA21x2_ASAP7_75t_R _4560_ (.A1(_0065_),
    .A2(net230),
    .B(_0064_),
    .Y(_1694_));
 OA21x2_ASAP7_75t_R _4561_ (.A1(_0042_),
    .A2(_1694_),
    .B(_0063_),
    .Y(_1695_));
 OA21x2_ASAP7_75t_R _4562_ (.A1(_0052_),
    .A2(_0059_),
    .B(_0058_),
    .Y(_1696_));
 OA21x2_ASAP7_75t_R _4563_ (.A1(_0746_),
    .A2(_1696_),
    .B(_0066_),
    .Y(_1697_));
 OA21x2_ASAP7_75t_R _4564_ (.A1(_1623_),
    .A2(_1697_),
    .B(_0079_),
    .Y(_1698_));
 OA21x2_ASAP7_75t_R _4565_ (.A1(_0744_),
    .A2(_1695_),
    .B(_1698_),
    .Y(_1699_));
 OA21x2_ASAP7_75t_R _4566_ (.A1(_0078_),
    .A2(net188),
    .B(_0077_),
    .Y(_1700_));
 OA21x2_ASAP7_75t_R _4567_ (.A1(_0032_),
    .A2(_1700_),
    .B(_0076_),
    .Y(_1701_));
 OA21x2_ASAP7_75t_R _4568_ (.A1(_0742_),
    .A2(_1701_),
    .B(_0075_),
    .Y(_1702_));
 OA21x2_ASAP7_75t_R _4569_ (.A1(_1637_),
    .A2(_1699_),
    .B(_1702_),
    .Y(_1703_));
 OA21x2_ASAP7_75t_R _4570_ (.A1(_0027_),
    .A2(_1703_),
    .B(_0074_),
    .Y(_1704_));
 OA21x2_ASAP7_75t_R _4571_ (.A1(net170),
    .A2(_1704_),
    .B(_0073_),
    .Y(_3554_));
 INVx2_ASAP7_75t_R _4572_ (.A(_1564_),
    .Y(_3189_));
 OA21x2_ASAP7_75t_R _4573_ (.A1(_0037_),
    .A2(_1699_),
    .B(_0078_),
    .Y(_1705_));
 OA21x2_ASAP7_75t_R _4574_ (.A1(net189),
    .A2(_1705_),
    .B(_0077_),
    .Y(_3193_));
 INVx2_ASAP7_75t_R _4575_ (.A(_1568_),
    .Y(_3517_));
 INVx2_ASAP7_75t_R _4576_ (.A(_1570_),
    .Y(_3519_));
 XNOR2x2_ASAP7_75t_R _4577_ (.A(_0085_),
    .B(net186),
    .Y(_1706_));
 OR2x2_ASAP7_75t_R _4578_ (.A(_1573_),
    .B(_1677_),
    .Y(_1707_));
 OA21x2_ASAP7_75t_R _4579_ (.A1(_1676_),
    .A2(_1706_),
    .B(_1707_),
    .Y(_3558_));
 INVx2_ASAP7_75t_R _4580_ (.A(_1575_),
    .Y(_3195_));
 AND2x2_ASAP7_75t_R _4581_ (.A(net39),
    .B(_1612_),
    .Y(_1708_));
 AND2x2_ASAP7_75t_R _4582_ (.A(_1508_),
    .B(_1614_),
    .Y(_1709_));
 OA21x2_ASAP7_75t_R _4583_ (.A1(_1708_),
    .A2(_1709_),
    .B(_3554_),
    .Y(_3575_));
 OR2x2_ASAP7_75t_R _4584_ (.A(_0017_),
    .B(_1620_),
    .Y(_1710_));
 NOR2x2_ASAP7_75t_R _4585_ (.A(_1508_),
    .B(_1710_),
    .Y(_1711_));
 AND3x2_ASAP7_75t_R _4586_ (.A(_1530_),
    .B(_1508_),
    .C(_1532_),
    .Y(_1712_));
 OR2x2_ASAP7_75t_R _4587_ (.A(_1544_),
    .B(net39),
    .Y(_1713_));
 OA211x2_ASAP7_75t_R _4588_ (.A1(_1508_),
    .A2(_1651_),
    .B(_3575_),
    .C(_1713_),
    .Y(_3573_));
 AND3x2_ASAP7_75t_R _4589_ (.A(_1652_),
    .B(net39),
    .C(_1671_),
    .Y(_1714_));
 AO21x2_ASAP7_75t_R _4590_ (.A1(_1542_),
    .A2(_1508_),
    .B(_1714_),
    .Y(_1715_));
 AND2x2_ASAP7_75t_R _4591_ (.A(_3573_),
    .B(_1715_),
    .Y(_3571_));
 AND2x2_ASAP7_75t_R _4592_ (.A(net39),
    .B(_1657_),
    .Y(_1716_));
 AO21x2_ASAP7_75t_R _4593_ (.A1(_1508_),
    .A2(_1537_),
    .B(_1716_),
    .Y(_1717_));
 AND2x2_ASAP7_75t_R _4594_ (.A(_3571_),
    .B(_1717_),
    .Y(_3569_));
 OA21x2_ASAP7_75t_R _4595_ (.A1(_1711_),
    .A2(_1712_),
    .B(_3569_),
    .Y(_3567_));
 AND2x2_ASAP7_75t_R _4596_ (.A(net39),
    .B(_1669_),
    .Y(_1718_));
 AO21x2_ASAP7_75t_R _4597_ (.A1(_1549_),
    .A2(_1508_),
    .B(_1718_),
    .Y(_1719_));
 AND2x2_ASAP7_75t_R _4598_ (.A(_3567_),
    .B(_1719_),
    .Y(_3563_));
 NOR3x2_ASAP7_75t_R _4599_ (.B(_1443_),
    .C(_1457_),
    .Y(_1720_),
    .A(_1432_));
 OA211x2_ASAP7_75t_R _4600_ (.A1(_1424_),
    .A2(_1498_),
    .B(_1534_),
    .C(_1535_),
    .Y(_1721_));
 AND5x2_ASAP7_75t_R _4601_ (.A(_1542_),
    .B(_1544_),
    .C(_1549_),
    .D(_1526_),
    .E(_1721_),
    .Y(_1722_));
 AND2x2_ASAP7_75t_R _4602_ (.A(_1720_),
    .B(_1722_),
    .Y(_1723_));
 OA21x2_ASAP7_75t_R _4603_ (.A1(_1723_),
    .A2(_1606_),
    .B(_3563_),
    .Y(_3561_));
 OA211x2_ASAP7_75t_R _4604_ (.A1(_1662_),
    .A2(_1665_),
    .B(_1667_),
    .C(_1507_),
    .Y(_1724_));
 AO21x2_ASAP7_75t_R _4605_ (.A1(_1553_),
    .A2(_1508_),
    .B(_1724_),
    .Y(_1725_));
 AND2x2_ASAP7_75t_R _4606_ (.A(_3567_),
    .B(_1725_),
    .Y(_3565_));
 INVx2_ASAP7_75t_R _4607_ (.A(_0108_),
    .Y(_1726_));
 AND2x2_ASAP7_75t_R _4608_ (.A(_1726_),
    .B(net38),
    .Y(_3576_));
 OR2x4_ASAP7_75t_R _4609_ (.A(_0110_),
    .B(net229),
    .Y(_1727_));
 TAPCELL_ASAP7_75t_R PHY_151 ();
 INVx2_ASAP7_75t_R _4611_ (.A(_1727_),
    .Y(_3579_));
 INVx2_ASAP7_75t_R _4612_ (.A(_0757_),
    .Y(_1728_));
 OA21x2_ASAP7_75t_R _4613_ (.A1(_1502_),
    .A2(_1503_),
    .B(_0762_),
    .Y(_1729_));
 INVx2_ASAP7_75t_R _4614_ (.A(_0762_),
    .Y(_1730_));
 AND3x2_ASAP7_75t_R _4615_ (.A(_1730_),
    .B(_1534_),
    .C(_1535_),
    .Y(_1731_));
 TAPCELL_ASAP7_75t_R PHY_150 ();
 INVx2_ASAP7_75t_R _4617_ (.A(_0764_),
    .Y(_1733_));
 OR2x2_ASAP7_75t_R _4618_ (.A(_1733_),
    .B(_0740_),
    .Y(_1734_));
 INVx2_ASAP7_75t_R _4619_ (.A(_0740_),
    .Y(_1735_));
 OR2x2_ASAP7_75t_R _4620_ (.A(_0764_),
    .B(_1735_),
    .Y(_1736_));
 AO221x2_ASAP7_75t_R _4621_ (.A1(_0488_),
    .A2(net162),
    .B1(_1734_),
    .B2(_1736_),
    .C(_1469_),
    .Y(_1737_));
 OR2x2_ASAP7_75t_R _4622_ (.A(_0764_),
    .B(_0740_),
    .Y(_1738_));
 NAND2x2_ASAP7_75t_R _4623_ (.A(_0764_),
    .B(_0740_),
    .Y(_1739_));
 AO221x2_ASAP7_75t_R _4624_ (.A1(_0488_),
    .A2(net162),
    .B1(_1738_),
    .B2(_1739_),
    .C(_1407_),
    .Y(_1740_));
 OR2x2_ASAP7_75t_R _4625_ (.A(_1469_),
    .B(_1738_),
    .Y(_1741_));
 OR2x2_ASAP7_75t_R _4626_ (.A(_1469_),
    .B(_1739_),
    .Y(_1742_));
 AO211x2_ASAP7_75t_R _4627_ (.A1(_1741_),
    .A2(_1742_),
    .B(_1646_),
    .C(net180),
    .Y(_1743_));
 OR3x2_ASAP7_75t_R _4628_ (.A(_1733_),
    .B(_0740_),
    .C(_1407_),
    .Y(_1744_));
 OR3x2_ASAP7_75t_R _4629_ (.A(_0764_),
    .B(_1735_),
    .C(_1407_),
    .Y(_1745_));
 AO211x2_ASAP7_75t_R _4630_ (.A1(_1744_),
    .A2(_1745_),
    .B(_1646_),
    .C(net180),
    .Y(_1746_));
 AND4x2_ASAP7_75t_R _4631_ (.A(_1737_),
    .B(_1740_),
    .C(_1743_),
    .D(_1746_),
    .Y(_1747_));
 OA211x2_ASAP7_75t_R _4632_ (.A1(_1729_),
    .A2(_1731_),
    .B(_1747_),
    .C(_1655_),
    .Y(_1748_));
 OR2x2_ASAP7_75t_R _4633_ (.A(_1733_),
    .B(_1469_),
    .Y(_1749_));
 OR2x2_ASAP7_75t_R _4634_ (.A(_0764_),
    .B(_1407_),
    .Y(_1750_));
 AO22x2_ASAP7_75t_R _4635_ (.A1(_0488_),
    .A2(net162),
    .B1(_1749_),
    .B2(_1750_),
    .Y(_1751_));
 OR4x2_ASAP7_75t_R _4636_ (.A(_1646_),
    .B(_0764_),
    .C(net209),
    .D(_1469_),
    .Y(_1752_));
 OR4x2_ASAP7_75t_R _4637_ (.A(_1646_),
    .B(_1733_),
    .C(net209),
    .D(_1407_),
    .Y(_1753_));
 AND3x2_ASAP7_75t_R _4638_ (.A(_1751_),
    .B(_1752_),
    .C(_1753_),
    .Y(_1754_));
 AO21x2_ASAP7_75t_R _4639_ (.A1(_1534_),
    .A2(_1535_),
    .B(_1730_),
    .Y(_1755_));
 OR3x2_ASAP7_75t_R _4640_ (.A(_0762_),
    .B(_1502_),
    .C(_1503_),
    .Y(_1756_));
 AND2x2_ASAP7_75t_R _4641_ (.A(_0738_),
    .B(_1735_),
    .Y(_1757_));
 AND4x2_ASAP7_75t_R _4642_ (.A(_1754_),
    .B(_1755_),
    .C(_1756_),
    .D(_1757_),
    .Y(_1758_));
 OR2x2_ASAP7_75t_R _4643_ (.A(_1748_),
    .B(_1758_),
    .Y(_1759_));
 AO221x2_ASAP7_75t_R _4644_ (.A1(_0738_),
    .A2(_0740_),
    .B1(_1720_),
    .B2(_1722_),
    .C(_1597_),
    .Y(_1760_));
 OR2x2_ASAP7_75t_R _4645_ (.A(_1729_),
    .B(_1731_),
    .Y(_1761_));
 NOR2x2_ASAP7_75t_R _4646_ (.A(_1754_),
    .B(_1761_),
    .Y(_1762_));
 AO32x2_ASAP7_75t_R _4647_ (.A1(_1506_),
    .A2(_1596_),
    .A3(_1759_),
    .B1(_1760_),
    .B2(_1762_),
    .Y(_1763_));
 AND2x2_ASAP7_75t_R _4648_ (.A(_0721_),
    .B(net162),
    .Y(_1764_));
 XOR2x2_ASAP7_75t_R _4649_ (.A(_0760_),
    .B(_1405_),
    .Y(_1765_));
 XNOR2x2_ASAP7_75t_R _4650_ (.A(_1764_),
    .B(_1765_),
    .Y(_1766_));
 XNOR2x2_ASAP7_75t_R _4651_ (.A(_0761_),
    .B(_1530_),
    .Y(_1767_));
 AO221x2_ASAP7_75t_R _4652_ (.A1(_0736_),
    .A2(_0737_),
    .B1(_1720_),
    .B2(_1722_),
    .C(_1597_),
    .Y(_1768_));
 XOR2x2_ASAP7_75t_R _4653_ (.A(_1764_),
    .B(_1765_),
    .Y(_1769_));
 INVx2_ASAP7_75t_R _4654_ (.A(_0761_),
    .Y(_1770_));
 OR2x2_ASAP7_75t_R _4655_ (.A(_1770_),
    .B(_0737_),
    .Y(_1771_));
 OR2x2_ASAP7_75t_R _4656_ (.A(_0761_),
    .B(_1619_),
    .Y(_1772_));
 AO22x2_ASAP7_75t_R _4657_ (.A1(_1528_),
    .A2(_1529_),
    .B1(_1771_),
    .B2(_1772_),
    .Y(_1773_));
 OR2x2_ASAP7_75t_R _4658_ (.A(_0761_),
    .B(_0737_),
    .Y(_1774_));
 OR2x2_ASAP7_75t_R _4659_ (.A(_1770_),
    .B(_1619_),
    .Y(_1775_));
 AO211x2_ASAP7_75t_R _4660_ (.A1(_1774_),
    .A2(_1775_),
    .B(_1441_),
    .C(_1442_),
    .Y(_1776_));
 NAND2x2_ASAP7_75t_R _4661_ (.A(_1773_),
    .B(_1776_),
    .Y(_1777_));
 AND3x2_ASAP7_75t_R _4662_ (.A(_0736_),
    .B(_1619_),
    .C(_1766_),
    .Y(_1778_));
 XNOR2x2_ASAP7_75t_R _4663_ (.A(_1770_),
    .B(_1530_),
    .Y(_1779_));
 AO32x2_ASAP7_75t_R _4664_ (.A1(_1663_),
    .A2(_1769_),
    .A3(_1777_),
    .B1(_1778_),
    .B2(_1779_),
    .Y(_1780_));
 AO32x2_ASAP7_75t_R _4665_ (.A1(_1766_),
    .A2(_1767_),
    .A3(_1768_),
    .B1(_1780_),
    .B2(net223),
    .Y(_1781_));
 XNOR2x2_ASAP7_75t_R _4666_ (.A(_0763_),
    .B(_1671_),
    .Y(_1782_));
 OA21x2_ASAP7_75t_R _4667_ (.A1(_1550_),
    .A2(_1551_),
    .B(_0758_),
    .Y(_1783_));
 INVx2_ASAP7_75t_R _4668_ (.A(_0758_),
    .Y(_1784_));
 AND3x2_ASAP7_75t_R _4669_ (.A(_1784_),
    .B(_1450_),
    .C(_1452_),
    .Y(_1785_));
 OA21x2_ASAP7_75t_R _4670_ (.A1(_1783_),
    .A2(_1785_),
    .B(_1602_),
    .Y(_1786_));
 INVx2_ASAP7_75t_R _4671_ (.A(_0021_),
    .Y(_1787_));
 INVx2_ASAP7_75t_R _4672_ (.A(_0754_),
    .Y(_1788_));
 AND2x2_ASAP7_75t_R _4673_ (.A(_1787_),
    .B(_1788_),
    .Y(_1789_));
 AND2x2_ASAP7_75t_R _4674_ (.A(_0021_),
    .B(_0754_),
    .Y(_1790_));
 OA21x2_ASAP7_75t_R _4675_ (.A1(_1789_),
    .A2(_1790_),
    .B(_1526_),
    .Y(_1791_));
 OR2x2_ASAP7_75t_R _4676_ (.A(_1547_),
    .B(_1548_),
    .Y(_1792_));
 AO33x2_ASAP7_75t_R _4677_ (.A1(_1659_),
    .A2(_0759_),
    .A3(_1792_),
    .B1(_1497_),
    .B2(_1788_),
    .B3(_0021_),
    .Y(_1793_));
 NOR3x2_ASAP7_75t_R _4678_ (.B(_1791_),
    .C(_1793_),
    .Y(_1794_),
    .A(_1786_));
 AO21x2_ASAP7_75t_R _4679_ (.A1(_1782_),
    .A2(_1794_),
    .B(net229),
    .Y(_1795_));
 OA22x2_ASAP7_75t_R _4680_ (.A1(_0763_),
    .A2(_1670_),
    .B1(_1497_),
    .B2(_0754_),
    .Y(_1796_));
 OR2x2_ASAP7_75t_R _4681_ (.A(net39),
    .B(_1796_),
    .Y(_1797_));
 INVx2_ASAP7_75t_R _4682_ (.A(_0759_),
    .Y(_1798_));
 AO22x2_ASAP7_75t_R _4683_ (.A1(_1784_),
    .A2(_1552_),
    .B1(_1792_),
    .B2(_1798_),
    .Y(_1799_));
 AND3x2_ASAP7_75t_R _4684_ (.A(_1720_),
    .B(_1722_),
    .C(_1799_),
    .Y(_1800_));
 OR2x2_ASAP7_75t_R _4685_ (.A(_0735_),
    .B(_1597_),
    .Y(_1801_));
 AND2x2_ASAP7_75t_R _4686_ (.A(_1480_),
    .B(_1482_),
    .Y(_1802_));
 XNOR2x2_ASAP7_75t_R _4687_ (.A(_0759_),
    .B(_1802_),
    .Y(_1803_));
 AND2x2_ASAP7_75t_R _4688_ (.A(_0763_),
    .B(_1597_),
    .Y(_1804_));
 AND2x2_ASAP7_75t_R _4689_ (.A(_1659_),
    .B(_1506_),
    .Y(_1805_));
 OA21x2_ASAP7_75t_R _4690_ (.A1(_0734_),
    .A2(_1597_),
    .B(_0758_),
    .Y(_1806_));
 AO32x2_ASAP7_75t_R _4691_ (.A1(_1798_),
    .A2(_1802_),
    .A3(_1805_),
    .B1(_1806_),
    .B2(_1600_),
    .Y(_1807_));
 AO221x2_ASAP7_75t_R _4692_ (.A1(_1801_),
    .A2(_1803_),
    .B1(_1804_),
    .B2(_1670_),
    .C(_1807_),
    .Y(_1808_));
 OR4x2_ASAP7_75t_R _4693_ (.A(_0084_),
    .B(_0087_),
    .C(_0756_),
    .D(_0755_),
    .Y(_1809_));
 OR5x2_ASAP7_75t_R _4694_ (.A(_0069_),
    .B(_0072_),
    .C(_0753_),
    .D(_0752_),
    .E(_1809_),
    .Y(_1810_));
 INVx2_ASAP7_75t_R _4695_ (.A(_0750_),
    .Y(_1811_));
 OA21x2_ASAP7_75t_R _4696_ (.A1(_0057_),
    .A2(_1811_),
    .B(_0107_),
    .Y(_1812_));
 OR2x2_ASAP7_75t_R _4697_ (.A(_0062_),
    .B(_0751_),
    .Y(_1813_));
 OA21x2_ASAP7_75t_R _4698_ (.A1(_0106_),
    .A2(_0751_),
    .B(_0105_),
    .Y(_1814_));
 OA21x2_ASAP7_75t_R _4699_ (.A1(_1812_),
    .A2(_1813_),
    .B(_1814_),
    .Y(_1815_));
 OA21x2_ASAP7_75t_R _4700_ (.A1(_0100_),
    .A2(_0756_),
    .B(_0099_),
    .Y(_1816_));
 OA21x2_ASAP7_75t_R _4701_ (.A1(_0084_),
    .A2(_1816_),
    .B(_0098_),
    .Y(_1817_));
 OA211x2_ASAP7_75t_R _4702_ (.A1(_0755_),
    .A2(_1817_),
    .B(_0096_),
    .C(_0097_),
    .Y(_1818_));
 OA21x2_ASAP7_75t_R _4703_ (.A1(_1810_),
    .A2(_1815_),
    .B(_1818_),
    .Y(_1819_));
 OA21x2_ASAP7_75t_R _4704_ (.A1(_0104_),
    .A2(_0753_),
    .B(_0103_),
    .Y(_1820_));
 OA21x2_ASAP7_75t_R _4705_ (.A1(_0069_),
    .A2(_1820_),
    .B(_0102_),
    .Y(_1821_));
 OA21x2_ASAP7_75t_R _4706_ (.A1(_0752_),
    .A2(_1821_),
    .B(_0101_),
    .Y(_1822_));
 OR2x2_ASAP7_75t_R _4707_ (.A(_1809_),
    .B(_1822_),
    .Y(_1823_));
 OR5x2_ASAP7_75t_R _4708_ (.A(_0057_),
    .B(_0055_),
    .C(_0083_),
    .D(_1810_),
    .E(_1813_),
    .Y(_1824_));
 INVx2_ASAP7_75t_R _4709_ (.A(_1824_),
    .Y(_1825_));
 AO221x2_ASAP7_75t_R _4710_ (.A1(_0083_),
    .A2(_0096_),
    .B1(_1819_),
    .B2(_1823_),
    .C(_1825_),
    .Y(_1826_));
 OA211x2_ASAP7_75t_R _4711_ (.A1(_0734_),
    .A2(_1597_),
    .B(_1552_),
    .C(_1784_),
    .Y(_1827_));
 OA211x2_ASAP7_75t_R _4712_ (.A1(_1787_),
    .A2(_1597_),
    .B(_1497_),
    .C(_0754_),
    .Y(_1828_));
 XOR2x2_ASAP7_75t_R _4713_ (.A(net171),
    .B(_0081_),
    .Y(_1829_));
 OR4x2_ASAP7_75t_R _4714_ (.A(_0080_),
    .B(_0090_),
    .C(_0091_),
    .D(_0092_),
    .Y(_1830_));
 OR3x2_ASAP7_75t_R _4715_ (.A(_0093_),
    .B(_0094_),
    .C(_1830_),
    .Y(_1831_));
 OR5x2_ASAP7_75t_R _4716_ (.A(_0088_),
    .B(_0089_),
    .C(_0095_),
    .D(_1829_),
    .E(_1831_),
    .Y(_1832_));
 OR4x2_ASAP7_75t_R _4717_ (.A(_1826_),
    .B(_1827_),
    .C(_1828_),
    .D(_1832_),
    .Y(_1833_));
 NOR3x2_ASAP7_75t_R _4718_ (.B(_1808_),
    .C(_1833_),
    .Y(_1834_),
    .A(_1800_));
 AND5x2_ASAP7_75t_R _4719_ (.A(_1763_),
    .B(_1781_),
    .C(_1795_),
    .D(_1797_),
    .E(_1834_),
    .Y(_1835_));
 OR2x2_ASAP7_75t_R _4720_ (.A(_1443_),
    .B(net39),
    .Y(_1836_));
 OR2x2_ASAP7_75t_R _4721_ (.A(_1508_),
    .B(_1621_),
    .Y(_1837_));
 OR2x2_ASAP7_75t_R _4722_ (.A(_1635_),
    .B(_1641_),
    .Y(_1838_));
 NAND2x2_ASAP7_75t_R _4723_ (.A(_1542_),
    .B(_1537_),
    .Y(_1839_));
 OR5x2_ASAP7_75t_R _4724_ (.A(_1472_),
    .B(_1491_),
    .C(net39),
    .D(_1838_),
    .E(_1839_),
    .Y(_1840_));
 OR3x2_ASAP7_75t_R _4725_ (.A(_0020_),
    .B(_1649_),
    .C(_1650_),
    .Y(_1841_));
 NAND2x2_ASAP7_75t_R _4726_ (.A(_1654_),
    .B(_1656_),
    .Y(_1842_));
 AO21x2_ASAP7_75t_R _4727_ (.A1(_1480_),
    .A2(_1482_),
    .B(_1659_),
    .Y(_1843_));
 OR3x2_ASAP7_75t_R _4728_ (.A(_0735_),
    .B(_1547_),
    .C(_1548_),
    .Y(_1844_));
 OA21x2_ASAP7_75t_R _4729_ (.A1(_1476_),
    .A2(net209),
    .B(_1664_),
    .Y(_1845_));
 AND3x2_ASAP7_75t_R _4730_ (.A(_0721_),
    .B(net162),
    .C(_1661_),
    .Y(_1846_));
 OR4x2_ASAP7_75t_R _4731_ (.A(_0015_),
    .B(_0016_),
    .C(_1845_),
    .D(_1846_),
    .Y(_1847_));
 AO21x2_ASAP7_75t_R _4732_ (.A1(_1843_),
    .A2(_1844_),
    .B(_1847_),
    .Y(_1848_));
 XNOR2x2_ASAP7_75t_R _4733_ (.A(_0739_),
    .B(_1670_),
    .Y(_1849_));
 OR5x2_ASAP7_75t_R _4734_ (.A(_0018_),
    .B(_0019_),
    .C(_1842_),
    .D(_1848_),
    .E(_1849_),
    .Y(_1850_));
 OR4x2_ASAP7_75t_R _4735_ (.A(net229),
    .B(_1838_),
    .C(_1841_),
    .D(_1850_),
    .Y(_1851_));
 OR3x2_ASAP7_75t_R _4736_ (.A(_0022_),
    .B(_1609_),
    .C(_1610_),
    .Y(_1852_));
 AO21x2_ASAP7_75t_R _4737_ (.A1(_1601_),
    .A2(_1605_),
    .B(_1852_),
    .Y(_1853_));
 OA22x2_ASAP7_75t_R _4738_ (.A1(net229),
    .A2(_1853_),
    .B1(_1615_),
    .B2(_1616_),
    .Y(_1854_));
 AO221x2_ASAP7_75t_R _4739_ (.A1(_1836_),
    .A2(_1837_),
    .B1(_1840_),
    .B2(_1851_),
    .C(_1854_),
    .Y(_1855_));
 TAPCELL_ASAP7_75t_R PHY_149 ();
 OA21x2_ASAP7_75t_R _4741_ (.A1(_1728_),
    .A2(_1835_),
    .B(_1855_),
    .Y(_1857_));
 XNOR2x2_ASAP7_75t_R _4742_ (.A(_0023_),
    .B(net168),
    .Y(_1858_));
 AND3x2_ASAP7_75t_R _4743_ (.A(net39),
    .B(_1858_),
    .C(_1612_),
    .Y(_1859_));
 AND3x2_ASAP7_75t_R _4744_ (.A(_3456_),
    .B(net229),
    .C(_1614_),
    .Y(_1860_));
 INVx2_ASAP7_75t_R _4745_ (.A(_1826_),
    .Y(_1861_));
 OA21x2_ASAP7_75t_R _4746_ (.A1(_1859_),
    .A2(_1860_),
    .B(_1861_),
    .Y(_1862_));
 AO21x2_ASAP7_75t_R _4747_ (.A1(_1674_),
    .A2(_1862_),
    .B(_1598_),
    .Y(_1863_));
 OR2x6_ASAP7_75t_R _4748_ (.A(_1857_),
    .B(_1863_),
    .Y(_1864_));
 TAPCELL_ASAP7_75t_R PHY_148 ();
 TAPCELL_ASAP7_75t_R PHY_147 ();
 TAPCELL_ASAP7_75t_R PHY_146 ();
 TAPCELL_ASAP7_75t_R PHY_145 ();
 AND2x2_ASAP7_75t_R _4753_ (.A(net38),
    .B(net222),
    .Y(_3209_));
 OA21x2_ASAP7_75t_R _4754_ (.A1(_0112_),
    .A2(_3208_),
    .B(_0111_),
    .Y(_1869_));
 OA21x2_ASAP7_75t_R _4755_ (.A1(_0765_),
    .A2(_1869_),
    .B(_0109_),
    .Y(_1870_));
 OR3x2_ASAP7_75t_R _4756_ (.A(_0552_),
    .B(_0553_),
    .C(_1870_),
    .Y(_1871_));
 OR3x2_ASAP7_75t_R _4757_ (.A(_0514_),
    .B(_0551_),
    .C(_1871_),
    .Y(_1872_));
 AO21x2_ASAP7_75t_R _4758_ (.A1(_0513_),
    .A2(_1872_),
    .B(_0512_),
    .Y(_1873_));
 AO21x2_ASAP7_75t_R _4759_ (.A1(_0511_),
    .A2(_1873_),
    .B(_0510_),
    .Y(_1874_));
 AND2x2_ASAP7_75t_R _4760_ (.A(_0509_),
    .B(_1874_),
    .Y(_3203_));
 OA21x2_ASAP7_75t_R _4761_ (.A1(_0508_),
    .A2(_3203_),
    .B(_0507_),
    .Y(_1875_));
 OA21x2_ASAP7_75t_R _4762_ (.A1(_0732_),
    .A2(_1875_),
    .B(_0506_),
    .Y(_3201_));
 OA21x2_ASAP7_75t_R _4763_ (.A1(_0505_),
    .A2(_3201_),
    .B(_0504_),
    .Y(_1876_));
 OA21x2_ASAP7_75t_R _4764_ (.A1(_0731_),
    .A2(_1876_),
    .B(_0503_),
    .Y(_3199_));
 INVx2_ASAP7_75t_R _4765_ (.A(_1871_),
    .Y(_3580_));
 CKINVDCx20_ASAP7_75t_R _4766_ (.A(_1864_),
    .Y(_1877_));
 TAPCELL_ASAP7_75t_R PHY_144 ();
 TAPCELL_ASAP7_75t_R PHY_143 ();
 AND2x2_ASAP7_75t_R _4769_ (.A(_0118_),
    .B(_1677_),
    .Y(_1879_));
 INVx2_ASAP7_75t_R _4770_ (.A(_0117_),
    .Y(_1880_));
 AND2x2_ASAP7_75t_R _4771_ (.A(_1880_),
    .B(net39),
    .Y(_1881_));
 AO21x2_ASAP7_75t_R _4772_ (.A1(_1207_),
    .A2(_1508_),
    .B(_1881_),
    .Y(_1882_));
 TAPCELL_ASAP7_75t_R PHY_142 ();
 NOR2x2_ASAP7_75t_R _4774_ (.A(_1677_),
    .B(_1882_),
    .Y(_1883_));
 OR3x2_ASAP7_75t_R _4775_ (.A(_1877_),
    .B(_1879_),
    .C(_1883_),
    .Y(_1884_));
 OA21x2_ASAP7_75t_R _4776_ (.A1(_0119_),
    .A2(_1864_),
    .B(_1884_),
    .Y(_3644_));
 OA21x2_ASAP7_75t_R _4777_ (.A1(_0135_),
    .A2(_3216_),
    .B(_0134_),
    .Y(_1885_));
 OA21x2_ASAP7_75t_R _4778_ (.A1(_0774_),
    .A2(_1885_),
    .B(_0133_),
    .Y(_3215_));
 OA21x2_ASAP7_75t_R _4779_ (.A1(_0132_),
    .A2(_3215_),
    .B(_0131_),
    .Y(_1886_));
 OA21x2_ASAP7_75t_R _4780_ (.A1(_0773_),
    .A2(_1886_),
    .B(_0130_),
    .Y(_3214_));
 OA21x2_ASAP7_75t_R _4781_ (.A1(_0129_),
    .A2(_3214_),
    .B(_0128_),
    .Y(_1887_));
 OA21x2_ASAP7_75t_R _4782_ (.A1(_0772_),
    .A2(_1887_),
    .B(_0127_),
    .Y(_3213_));
 OA21x2_ASAP7_75t_R _4783_ (.A1(_0126_),
    .A2(_3213_),
    .B(_0125_),
    .Y(_1888_));
 OA21x2_ASAP7_75t_R _4784_ (.A1(_0771_),
    .A2(_1888_),
    .B(_0124_),
    .Y(_3211_));
 OA21x2_ASAP7_75t_R _4785_ (.A1(_0123_),
    .A2(_3211_),
    .B(_0122_),
    .Y(_1889_));
 OR2x2_ASAP7_75t_R _4786_ (.A(_0770_),
    .B(_1889_),
    .Y(_1890_));
 NAND2x2_ASAP7_75t_R _4787_ (.A(_0121_),
    .B(_1890_),
    .Y(_3588_));
 AND3x2_ASAP7_75t_R _4788_ (.A(_1348_),
    .B(_3239_),
    .C(_3588_),
    .Y(_3586_));
 INVx2_ASAP7_75t_R _4789_ (.A(_0137_),
    .Y(_1891_));
 AND2x2_ASAP7_75t_R _4790_ (.A(_1891_),
    .B(net38),
    .Y(_3599_));
 XNOR2x2_ASAP7_75t_R _4791_ (.A(_0776_),
    .B(_1348_),
    .Y(_1892_));
 NAND2x2_ASAP7_75t_R _4792_ (.A(net223),
    .B(_1892_),
    .Y(_1893_));
 INVx2_ASAP7_75t_R _4793_ (.A(_1893_),
    .Y(_3587_));
 INVx2_ASAP7_75t_R _4794_ (.A(_0139_),
    .Y(_1894_));
 AND2x2_ASAP7_75t_R _4795_ (.A(_1894_),
    .B(net223),
    .Y(_3221_));
 AND2x2_ASAP7_75t_R _4796_ (.A(_0586_),
    .B(net38),
    .Y(_1895_));
 AND2x2_ASAP7_75t_R _4797_ (.A(_1348_),
    .B(net229),
    .Y(_1896_));
 OR2x2_ASAP7_75t_R _4798_ (.A(_1895_),
    .B(_1896_),
    .Y(_1897_));
 TAPCELL_ASAP7_75t_R PHY_141 ();
 INVx2_ASAP7_75t_R _4800_ (.A(_1897_),
    .Y(_3223_));
 NOR2x2_ASAP7_75t_R _4801_ (.A(_1363_),
    .B(net38),
    .Y(_1898_));
 AO21x2_ASAP7_75t_R _4802_ (.A1(_0588_),
    .A2(net38),
    .B(_1898_),
    .Y(_1899_));
 TAPCELL_ASAP7_75t_R PHY_140 ();
 INVx2_ASAP7_75t_R _4804_ (.A(_1899_),
    .Y(_3225_));
 OR2x2_ASAP7_75t_R _4805_ (.A(_0590_),
    .B(_1508_),
    .Y(_1900_));
 OA21x2_ASAP7_75t_R _4806_ (.A1(_1388_),
    .A2(net38),
    .B(_1900_),
    .Y(_1901_));
 TAPCELL_ASAP7_75t_R PHY_139 ();
 INVx2_ASAP7_75t_R _4808_ (.A(_1901_),
    .Y(_3227_));
 AND2x2_ASAP7_75t_R _4809_ (.A(_0592_),
    .B(net39),
    .Y(_1902_));
 OA211x2_ASAP7_75t_R _4810_ (.A1(_1239_),
    .A2(_1248_),
    .B(_1508_),
    .C(_1257_),
    .Y(_1903_));
 OR2x2_ASAP7_75t_R _4811_ (.A(_1902_),
    .B(_1903_),
    .Y(_1904_));
 TAPCELL_ASAP7_75t_R PHY_138 ();
 INVx2_ASAP7_75t_R _4813_ (.A(_1904_),
    .Y(_3229_));
 OA211x2_ASAP7_75t_R _4814_ (.A1(_1458_),
    .A2(_1505_),
    .B(_0594_),
    .C(_1506_),
    .Y(_1905_));
 AO21x2_ASAP7_75t_R _4815_ (.A1(_1314_),
    .A2(_1508_),
    .B(_1905_),
    .Y(_1906_));
 TAPCELL_ASAP7_75t_R PHY_137 ();
 INVx2_ASAP7_75t_R _4817_ (.A(_1906_),
    .Y(_3231_));
 OA21x2_ASAP7_75t_R _4818_ (.A1(_0156_),
    .A2(_3232_),
    .B(_0155_),
    .Y(_1907_));
 OA21x2_ASAP7_75t_R _4819_ (.A1(_0781_),
    .A2(_1907_),
    .B(_0154_),
    .Y(_3230_));
 OA21x2_ASAP7_75t_R _4820_ (.A1(_0153_),
    .A2(_3230_),
    .B(_0152_),
    .Y(_1908_));
 OA21x2_ASAP7_75t_R _4821_ (.A1(_0780_),
    .A2(_1908_),
    .B(_0151_),
    .Y(_3228_));
 OA21x2_ASAP7_75t_R _4822_ (.A1(_0150_),
    .A2(_3228_),
    .B(_0149_),
    .Y(_1909_));
 OA21x2_ASAP7_75t_R _4823_ (.A1(_0779_),
    .A2(_1909_),
    .B(_0148_),
    .Y(_3226_));
 TAPCELL_ASAP7_75t_R PHY_136 ();
 TAPCELL_ASAP7_75t_R PHY_135 ();
 OR3x2_ASAP7_75t_R _4826_ (.A(_0147_),
    .B(_0778_),
    .C(_0779_),
    .Y(_1912_));
 OR2x2_ASAP7_75t_R _4827_ (.A(_0147_),
    .B(_0148_),
    .Y(_1913_));
 AO21x2_ASAP7_75t_R _4828_ (.A1(_0146_),
    .A2(_1913_),
    .B(_0778_),
    .Y(_1914_));
 AND3x2_ASAP7_75t_R _4829_ (.A(_0143_),
    .B(_0142_),
    .C(_0145_),
    .Y(_1915_));
 OA211x2_ASAP7_75t_R _4830_ (.A1(_1909_),
    .A2(_1912_),
    .B(_1914_),
    .C(_1915_),
    .Y(_1916_));
 AND3x2_ASAP7_75t_R _4831_ (.A(_0143_),
    .B(_0142_),
    .C(_0144_),
    .Y(_1917_));
 AO21x2_ASAP7_75t_R _4832_ (.A1(_0142_),
    .A2(_0777_),
    .B(_1917_),
    .Y(_1918_));
 OR4x2_ASAP7_75t_R _4833_ (.A(_0141_),
    .B(_0775_),
    .C(_1916_),
    .D(_1918_),
    .Y(_1919_));
 OA21x2_ASAP7_75t_R _4834_ (.A1(_0140_),
    .A2(_0775_),
    .B(_0138_),
    .Y(_1920_));
 AND2x2_ASAP7_75t_R _4835_ (.A(_1919_),
    .B(_1920_),
    .Y(_1921_));
 OR3x2_ASAP7_75t_R _4836_ (.A(_0136_),
    .B(_0137_),
    .C(net229),
    .Y(_1922_));
 OR4x2_ASAP7_75t_R _4837_ (.A(_1598_),
    .B(net234),
    .C(_1921_),
    .D(_1922_),
    .Y(_1923_));
 INVx2_ASAP7_75t_R _4838_ (.A(_1923_),
    .Y(_3609_));
 OR2x2_ASAP7_75t_R _4839_ (.A(_0158_),
    .B(net219),
    .Y(_1924_));
 OR3x2_ASAP7_75t_R _4840_ (.A(_0137_),
    .B(net229),
    .C(_1677_),
    .Y(_1925_));
 NAND2x2_ASAP7_75t_R _4841_ (.A(_1924_),
    .B(_1925_),
    .Y(_3611_));
 INVx2_ASAP7_75t_R _4842_ (.A(_0160_),
    .Y(_1926_));
 OA21x2_ASAP7_75t_R _4843_ (.A1(_0733_),
    .A2(_1723_),
    .B(_1506_),
    .Y(_1927_));
 TAPCELL_ASAP7_75t_R PHY_134 ();
 TAPCELL_ASAP7_75t_R PHY_133 ();
 AND3x2_ASAP7_75t_R _4846_ (.A(_1926_),
    .B(_1927_),
    .C(_1855_),
    .Y(_1930_));
 OA21x2_ASAP7_75t_R _4847_ (.A1(_1598_),
    .A2(_1674_),
    .B(_3221_),
    .Y(_1931_));
 OR2x2_ASAP7_75t_R _4848_ (.A(_1930_),
    .B(_1931_),
    .Y(_1932_));
 TAPCELL_ASAP7_75t_R PHY_132 ();
 INVx2_ASAP7_75t_R _4850_ (.A(_1932_),
    .Y(_3236_));
 OA211x2_ASAP7_75t_R _4851_ (.A1(_1909_),
    .A2(_1912_),
    .B(_1914_),
    .C(_0145_),
    .Y(_3224_));
 INVx2_ASAP7_75t_R _4852_ (.A(_0598_),
    .Y(_1933_));
 AND2x2_ASAP7_75t_R _4853_ (.A(net219),
    .B(_3225_),
    .Y(_1934_));
 AO21x2_ASAP7_75t_R _4854_ (.A1(_1933_),
    .A2(_1677_),
    .B(_1934_),
    .Y(_1935_));
 TAPCELL_ASAP7_75t_R PHY_131 ();
 OR2x2_ASAP7_75t_R _4856_ (.A(_1677_),
    .B(_1904_),
    .Y(_1936_));
 OA21x2_ASAP7_75t_R _4857_ (.A1(_0602_),
    .A2(net219),
    .B(_1936_),
    .Y(_3606_));
 INVx2_ASAP7_75t_R _4858_ (.A(_3606_),
    .Y(_3247_));
 OR2x2_ASAP7_75t_R _4859_ (.A(_1677_),
    .B(_1906_),
    .Y(_1937_));
 OA21x2_ASAP7_75t_R _4860_ (.A1(_0604_),
    .A2(net221),
    .B(_1937_),
    .Y(_3608_));
 INVx2_ASAP7_75t_R _4861_ (.A(_3608_),
    .Y(_3249_));
 OA21x2_ASAP7_75t_R _4862_ (.A1(_0177_),
    .A2(_3250_),
    .B(_0176_),
    .Y(_1938_));
 OA21x2_ASAP7_75t_R _4863_ (.A1(_0787_),
    .A2(_1938_),
    .B(_0175_),
    .Y(_3248_));
 OA21x2_ASAP7_75t_R _4864_ (.A1(_0174_),
    .A2(_3248_),
    .B(_0173_),
    .Y(_1939_));
 OA21x2_ASAP7_75t_R _4865_ (.A1(_0786_),
    .A2(_1939_),
    .B(_0172_),
    .Y(_1940_));
 OA21x2_ASAP7_75t_R _4866_ (.A1(_0171_),
    .A2(_1940_),
    .B(_0170_),
    .Y(_1941_));
 OA21x2_ASAP7_75t_R _4867_ (.A1(_0785_),
    .A2(_1941_),
    .B(_0169_),
    .Y(_3243_));
 NOR2x2_ASAP7_75t_R _4868_ (.A(_1748_),
    .B(_1758_),
    .Y(_1942_));
 OA221x2_ASAP7_75t_R _4869_ (.A1(_1655_),
    .A2(_1735_),
    .B1(_1458_),
    .B2(_1505_),
    .C(_1506_),
    .Y(_1943_));
 OA33x2_ASAP7_75t_R _4870_ (.A1(_1597_),
    .A2(_1723_),
    .A3(_1942_),
    .B1(_1943_),
    .B2(_1754_),
    .B3(_1761_),
    .Y(_1944_));
 OR3x2_ASAP7_75t_R _4871_ (.A(_1663_),
    .B(_0737_),
    .C(_1769_),
    .Y(_1945_));
 AO21x2_ASAP7_75t_R _4872_ (.A1(_1773_),
    .A2(_1776_),
    .B(_0736_),
    .Y(_1946_));
 OA22x2_ASAP7_75t_R _4873_ (.A1(_1767_),
    .A2(_1945_),
    .B1(_1946_),
    .B2(_1766_),
    .Y(_1947_));
 OA221x2_ASAP7_75t_R _4874_ (.A1(_1663_),
    .A2(_1619_),
    .B1(_1458_),
    .B2(_1505_),
    .C(_1506_),
    .Y(_1948_));
 OA33x2_ASAP7_75t_R _4875_ (.A1(_1597_),
    .A2(_1723_),
    .A3(_1947_),
    .B1(_1948_),
    .B2(_1769_),
    .B3(_1779_),
    .Y(_1949_));
 XNOR2x2_ASAP7_75t_R _4876_ (.A(_0763_),
    .B(_1849_),
    .Y(_1950_));
 OR3x2_ASAP7_75t_R _4877_ (.A(_1786_),
    .B(_1791_),
    .C(_1793_),
    .Y(_1951_));
 OA21x2_ASAP7_75t_R _4878_ (.A1(_1950_),
    .A2(_1951_),
    .B(net39),
    .Y(_1952_));
 NOR2x2_ASAP7_75t_R _4879_ (.A(net39),
    .B(_1796_),
    .Y(_1953_));
 OR3x2_ASAP7_75t_R _4880_ (.A(_1800_),
    .B(_1808_),
    .C(_1833_),
    .Y(_1954_));
 OR5x2_ASAP7_75t_R _4881_ (.A(_1944_),
    .B(_1949_),
    .C(_1952_),
    .D(_1953_),
    .E(_1954_),
    .Y(_1955_));
 AO21x2_ASAP7_75t_R _4882_ (.A1(_0757_),
    .A2(_1955_),
    .B(net234),
    .Y(_1956_));
 TAPCELL_ASAP7_75t_R PHY_130 ();
 OR3x2_ASAP7_75t_R _4884_ (.A(net229),
    .B(_1560_),
    .C(_1852_),
    .Y(_1958_));
 OR3x2_ASAP7_75t_R _4885_ (.A(_3457_),
    .B(net39),
    .C(_1615_),
    .Y(_1959_));
 AO21x2_ASAP7_75t_R _4886_ (.A1(_1958_),
    .A2(_1959_),
    .B(_1826_),
    .Y(_1960_));
 OA21x2_ASAP7_75t_R _4887_ (.A1(_1855_),
    .A2(_1960_),
    .B(_1927_),
    .Y(_1961_));
 TAPCELL_ASAP7_75t_R PHY_129 ();
 AO21x2_ASAP7_75t_R _4889_ (.A1(_1956_),
    .A2(_1961_),
    .B(_1923_),
    .Y(_1963_));
 OA21x2_ASAP7_75t_R _4890_ (.A1(_0180_),
    .A2(net222),
    .B(_1963_),
    .Y(_3614_));
 OA21x2_ASAP7_75t_R _4891_ (.A1(_0168_),
    .A2(_3243_),
    .B(_0167_),
    .Y(_1964_));
 OA21x2_ASAP7_75t_R _4892_ (.A1(_0784_),
    .A2(_1964_),
    .B(_0166_),
    .Y(_1965_));
 OA21x2_ASAP7_75t_R _4893_ (.A1(_0165_),
    .A2(_1965_),
    .B(_0164_),
    .Y(_1966_));
 OA21x2_ASAP7_75t_R _4894_ (.A1(_0783_),
    .A2(_1966_),
    .B(_0163_),
    .Y(_3237_));
 XNOR2x2_ASAP7_75t_R _4895_ (.A(_0770_),
    .B(_0585_),
    .Y(_1967_));
 AND2x2_ASAP7_75t_R _4896_ (.A(net38),
    .B(_1967_),
    .Y(_1968_));
 AO21x2_ASAP7_75t_R _4897_ (.A1(_3154_),
    .A2(net229),
    .B(_1968_),
    .Y(_3589_));
 AO21x2_ASAP7_75t_R _4898_ (.A1(_1927_),
    .A2(_1855_),
    .B(_3589_),
    .Y(_1969_));
 XNOR2x2_ASAP7_75t_R _4899_ (.A(_0595_),
    .B(_0777_),
    .Y(_1970_));
 OR3x2_ASAP7_75t_R _4900_ (.A(_1598_),
    .B(_1674_),
    .C(_1970_),
    .Y(_1971_));
 NAND2x2_ASAP7_75t_R _4901_ (.A(_1969_),
    .B(_1971_),
    .Y(_1972_));
 INVx2_ASAP7_75t_R _4902_ (.A(_1972_),
    .Y(_3601_));
 OR3x2_ASAP7_75t_R _4903_ (.A(_0596_),
    .B(_1598_),
    .C(_1674_),
    .Y(_1973_));
 AO21x2_ASAP7_75t_R _4904_ (.A1(_1927_),
    .A2(_1855_),
    .B(_1897_),
    .Y(_1974_));
 NAND2x2_ASAP7_75t_R _4905_ (.A(_1973_),
    .B(_1974_),
    .Y(_1975_));
 INVx2_ASAP7_75t_R _4906_ (.A(_1975_),
    .Y(_3240_));
 XNOR2x2_ASAP7_75t_R _4907_ (.A(_0597_),
    .B(_0778_),
    .Y(_1976_));
 XNOR2x2_ASAP7_75t_R _4908_ (.A(_0771_),
    .B(_0587_),
    .Y(_1977_));
 AND2x2_ASAP7_75t_R _4909_ (.A(net38),
    .B(_1977_),
    .Y(_1978_));
 AO21x2_ASAP7_75t_R _4910_ (.A1(_3239_),
    .A2(net229),
    .B(_1978_),
    .Y(_3591_));
 AND2x2_ASAP7_75t_R _4911_ (.A(net219),
    .B(_3591_),
    .Y(_1979_));
 AO21x2_ASAP7_75t_R _4912_ (.A1(_1677_),
    .A2(_1976_),
    .B(_1979_),
    .Y(_1980_));
 TAPCELL_ASAP7_75t_R PHY_128 ();
 INVx2_ASAP7_75t_R _4914_ (.A(_1935_),
    .Y(_3603_));
 XNOR2x2_ASAP7_75t_R _4915_ (.A(_0599_),
    .B(_0779_),
    .Y(_1981_));
 OR2x2_ASAP7_75t_R _4916_ (.A(_3159_),
    .B(net38),
    .Y(_1982_));
 XOR2x2_ASAP7_75t_R _4917_ (.A(_0589_),
    .B(_0772_),
    .Y(_1983_));
 OR2x2_ASAP7_75t_R _4918_ (.A(_1508_),
    .B(_1983_),
    .Y(_1984_));
 NAND2x2_ASAP7_75t_R _4919_ (.A(_1982_),
    .B(_1984_),
    .Y(_3593_));
 AND2x2_ASAP7_75t_R _4920_ (.A(net219),
    .B(_3593_),
    .Y(_1985_));
 AO21x2_ASAP7_75t_R _4921_ (.A1(_1677_),
    .A2(_1981_),
    .B(_1985_),
    .Y(_1986_));
 TAPCELL_ASAP7_75t_R PHY_127 ();
 AND2x2_ASAP7_75t_R _4923_ (.A(net219),
    .B(_1901_),
    .Y(_1987_));
 AO21x2_ASAP7_75t_R _4924_ (.A1(_0600_),
    .A2(_1677_),
    .B(_1987_),
    .Y(_3245_));
 AND2x2_ASAP7_75t_R _4925_ (.A(_3244_),
    .B(_1508_),
    .Y(_1988_));
 XNOR2x2_ASAP7_75t_R _4926_ (.A(_0773_),
    .B(_0591_),
    .Y(_1989_));
 AND2x2_ASAP7_75t_R _4927_ (.A(net39),
    .B(_1989_),
    .Y(_1990_));
 NOR2x2_ASAP7_75t_R _4928_ (.A(_1988_),
    .B(_1990_),
    .Y(_1991_));
 INVx2_ASAP7_75t_R _4929_ (.A(_1991_),
    .Y(_3595_));
 XOR2x2_ASAP7_75t_R _4930_ (.A(_0601_),
    .B(_0780_),
    .Y(_1992_));
 AND2x2_ASAP7_75t_R _4931_ (.A(_1927_),
    .B(_1992_),
    .Y(_1993_));
 NAND2x2_ASAP7_75t_R _4932_ (.A(_1855_),
    .B(_1993_),
    .Y(_1994_));
 OA21x2_ASAP7_75t_R _4933_ (.A1(_1677_),
    .A2(_3595_),
    .B(_1994_),
    .Y(_3605_));
 INVx2_ASAP7_75t_R _4934_ (.A(_0157_),
    .Y(_1995_));
 AND2x2_ASAP7_75t_R _4935_ (.A(_1995_),
    .B(net39),
    .Y(_1996_));
 AO21x2_ASAP7_75t_R _4936_ (.A1(_1336_),
    .A2(_1508_),
    .B(_1996_),
    .Y(_3234_));
 INVx2_ASAP7_75t_R _4937_ (.A(_0178_),
    .Y(_1997_));
 OR2x2_ASAP7_75t_R _4938_ (.A(_1997_),
    .B(net221),
    .Y(_1998_));
 OA21x2_ASAP7_75t_R _4939_ (.A1(_1677_),
    .A2(_3234_),
    .B(_1998_),
    .Y(_3252_));
 INVx2_ASAP7_75t_R _4940_ (.A(_0188_),
    .Y(_1999_));
 TAPCELL_ASAP7_75t_R PHY_126 ();
 AND2x2_ASAP7_75t_R _4942_ (.A(_1999_),
    .B(_1877_),
    .Y(_2001_));
 AO21x2_ASAP7_75t_R _4943_ (.A1(_1864_),
    .A2(_3252_),
    .B(_2001_),
    .Y(_2002_));
 INVx2_ASAP7_75t_R _4944_ (.A(_2002_),
    .Y(_3645_));
 INVx2_ASAP7_75t_R _4945_ (.A(_0811_),
    .Y(_3642_));
 TAPCELL_ASAP7_75t_R PHY_125 ();
 TAPCELL_ASAP7_75t_R PHY_124 ();
 XNOR2x2_ASAP7_75t_R _4948_ (.A(_0159_),
    .B(_0775_),
    .Y(_2005_));
 OR2x2_ASAP7_75t_R _4949_ (.A(_0605_),
    .B(_2005_),
    .Y(_2006_));
 INVx2_ASAP7_75t_R _4950_ (.A(_0605_),
    .Y(_2007_));
 XOR2x2_ASAP7_75t_R _4951_ (.A(_0159_),
    .B(_0775_),
    .Y(_2008_));
 OR2x2_ASAP7_75t_R _4952_ (.A(_2007_),
    .B(_2008_),
    .Y(_2009_));
 AO211x2_ASAP7_75t_R _4953_ (.A1(_2006_),
    .A2(_2009_),
    .B(_1598_),
    .C(net226),
    .Y(_2010_));
 OR2x2_ASAP7_75t_R _4954_ (.A(_2007_),
    .B(_3587_),
    .Y(_2011_));
 OR2x2_ASAP7_75t_R _4955_ (.A(_0605_),
    .B(_1893_),
    .Y(_2012_));
 AO22x2_ASAP7_75t_R _4956_ (.A1(_1927_),
    .A2(_1855_),
    .B1(_2011_),
    .B2(_2012_),
    .Y(_2013_));
 NAND3x2_ASAP7_75t_R _4957_ (.B(_2010_),
    .C(_2013_),
    .Y(_2014_),
    .A(_0606_));
 AO221x2_ASAP7_75t_R _4958_ (.A1(_1926_),
    .A2(_1677_),
    .B1(_1956_),
    .B2(_1961_),
    .C(_1931_),
    .Y(_2015_));
 OA21x2_ASAP7_75t_R _4959_ (.A1(_1598_),
    .A2(net226),
    .B(_3587_),
    .Y(_2016_));
 AO21x2_ASAP7_75t_R _4960_ (.A1(_1677_),
    .A2(_2008_),
    .B(_2016_),
    .Y(_2017_));
 OA22x2_ASAP7_75t_R _4961_ (.A1(net228),
    .A2(_2014_),
    .B1(_2015_),
    .B2(_2017_),
    .Y(_2018_));
 AND2x2_ASAP7_75t_R _4962_ (.A(_0757_),
    .B(_1955_),
    .Y(_2019_));
 OA22x2_ASAP7_75t_R _4963_ (.A1(_2019_),
    .A2(_1994_),
    .B1(_3595_),
    .B2(_1961_),
    .Y(_2020_));
 OA211x2_ASAP7_75t_R _4964_ (.A1(_1272_),
    .A2(_1289_),
    .B(_1508_),
    .C(_1291_),
    .Y(_2021_));
 XNOR2x2_ASAP7_75t_R _4965_ (.A(_0593_),
    .B(_0774_),
    .Y(_2022_));
 AND2x2_ASAP7_75t_R _4966_ (.A(net39),
    .B(_2022_),
    .Y(_2023_));
 OR4x2_ASAP7_75t_R _4967_ (.A(_0811_),
    .B(_1906_),
    .C(_2021_),
    .D(_2023_),
    .Y(_2024_));
 AO21x2_ASAP7_75t_R _4968_ (.A1(_1927_),
    .A2(_1855_),
    .B(_2024_),
    .Y(_2025_));
 XNOR2x2_ASAP7_75t_R _4969_ (.A(_0603_),
    .B(_0781_),
    .Y(_2026_));
 OR5x2_ASAP7_75t_R _4970_ (.A(_0811_),
    .B(_0604_),
    .C(_1598_),
    .D(net234),
    .E(_2026_),
    .Y(_2027_));
 AND2x2_ASAP7_75t_R _4971_ (.A(_2025_),
    .B(_2027_),
    .Y(_2028_));
 OR3x2_ASAP7_75t_R _4972_ (.A(_1901_),
    .B(_1904_),
    .C(_3593_),
    .Y(_2029_));
 OR3x2_ASAP7_75t_R _4973_ (.A(_0602_),
    .B(_0600_),
    .C(_1981_),
    .Y(_2030_));
 OR3x2_ASAP7_75t_R _4974_ (.A(_1598_),
    .B(net226),
    .C(_2030_),
    .Y(_2031_));
 OA21x2_ASAP7_75t_R _4975_ (.A1(_1677_),
    .A2(_2029_),
    .B(_2031_),
    .Y(_2032_));
 XNOR2x2_ASAP7_75t_R _4976_ (.A(_0787_),
    .B(_0609_),
    .Y(_2033_));
 XNOR2x2_ASAP7_75t_R _4977_ (.A(_0608_),
    .B(_0786_),
    .Y(_2034_));
 OR4x2_ASAP7_75t_R _4978_ (.A(_0187_),
    .B(_0811_),
    .C(_2033_),
    .D(_2034_),
    .Y(_2035_));
 XOR2x2_ASAP7_75t_R _4979_ (.A(_0184_),
    .B(_0785_),
    .Y(_2036_));
 OR3x2_ASAP7_75t_R _4980_ (.A(_0185_),
    .B(_0186_),
    .C(_2036_),
    .Y(_2037_));
 OR4x2_ASAP7_75t_R _4981_ (.A(_1857_),
    .B(_1863_),
    .C(_2035_),
    .D(_2037_),
    .Y(_2038_));
 OA31x2_ASAP7_75t_R _4982_ (.A1(_2020_),
    .A2(_2028_),
    .A3(_2032_),
    .B1(_2038_),
    .Y(_2039_));
 OR4x2_ASAP7_75t_R _4983_ (.A(_0598_),
    .B(_1598_),
    .C(net226),
    .D(_1976_),
    .Y(_2040_));
 AO211x2_ASAP7_75t_R _4984_ (.A1(_1927_),
    .A2(_1855_),
    .B(_1899_),
    .C(_3591_),
    .Y(_2041_));
 AO22x2_ASAP7_75t_R _4985_ (.A1(_1956_),
    .A2(_1961_),
    .B1(_2040_),
    .B2(_2041_),
    .Y(_2042_));
 INVx2_ASAP7_75t_R _4986_ (.A(_0183_),
    .Y(_2043_));
 XOR2x2_ASAP7_75t_R _4987_ (.A(_0607_),
    .B(_0784_),
    .Y(_2044_));
 NAND2x2_ASAP7_75t_R _4988_ (.A(_2043_),
    .B(_2044_),
    .Y(_2045_));
 OR3x2_ASAP7_75t_R _4989_ (.A(_1857_),
    .B(_1863_),
    .C(_2045_),
    .Y(_2046_));
 AND2x2_ASAP7_75t_R _4990_ (.A(_2042_),
    .B(_2046_),
    .Y(_2047_));
 INVx2_ASAP7_75t_R _4991_ (.A(_0182_),
    .Y(_2048_));
 XNOR2x2_ASAP7_75t_R _4992_ (.A(_0181_),
    .B(_0783_),
    .Y(_2049_));
 NAND2x2_ASAP7_75t_R _4993_ (.A(_2048_),
    .B(_2049_),
    .Y(_2050_));
 AO22x2_ASAP7_75t_R _4994_ (.A1(_1956_),
    .A2(_1961_),
    .B1(_1969_),
    .B2(_1971_),
    .Y(_2051_));
 OA22x2_ASAP7_75t_R _4995_ (.A1(net228),
    .A2(_2050_),
    .B1(_2051_),
    .B2(_3240_),
    .Y(_2052_));
 OR4x2_ASAP7_75t_R _4996_ (.A(_2018_),
    .B(_2039_),
    .C(_2047_),
    .D(_2052_),
    .Y(_2053_));
 AND3x2_ASAP7_75t_R _4997_ (.A(_0789_),
    .B(_1956_),
    .C(_1961_),
    .Y(_2054_));
 AO31x2_ASAP7_75t_R _4998_ (.A1(net228),
    .A2(_1924_),
    .A3(_1925_),
    .B(_2054_),
    .Y(_2055_));
 TAPCELL_ASAP7_75t_R PHY_123 ();
 OR2x2_ASAP7_75t_R _5000_ (.A(_1728_),
    .B(_1835_),
    .Y(_2056_));
 AO221x2_ASAP7_75t_R _5001_ (.A1(_0179_),
    .A2(_0180_),
    .B1(_1855_),
    .B2(_2056_),
    .C(_1863_),
    .Y(_2057_));
 INVx2_ASAP7_75t_R _5002_ (.A(_0788_),
    .Y(_2058_));
 INVx2_ASAP7_75t_R _5003_ (.A(_0782_),
    .Y(_2059_));
 OR2x2_ASAP7_75t_R _5004_ (.A(_0136_),
    .B(net229),
    .Y(_2060_));
 AO31x2_ASAP7_75t_R _5005_ (.A1(_2059_),
    .A2(_1927_),
    .A3(_1855_),
    .B(_2060_),
    .Y(_2061_));
 INVx2_ASAP7_75t_R _5006_ (.A(_0136_),
    .Y(_2062_));
 AND2x2_ASAP7_75t_R _5007_ (.A(_2062_),
    .B(net38),
    .Y(_2063_));
 OR4x2_ASAP7_75t_R _5008_ (.A(_0782_),
    .B(_1598_),
    .C(net226),
    .D(_2063_),
    .Y(_2064_));
 AO32x2_ASAP7_75t_R _5009_ (.A1(_2058_),
    .A2(_1956_),
    .A3(_1961_),
    .B1(_2061_),
    .B2(_2064_),
    .Y(_2065_));
 TAPCELL_ASAP7_75t_R PHY_122 ();
 OA31x2_ASAP7_75t_R _5011_ (.A1(_0782_),
    .A2(_1598_),
    .A3(net234),
    .B1(_2063_),
    .Y(_2067_));
 AND4x2_ASAP7_75t_R _5012_ (.A(_2059_),
    .B(_1927_),
    .C(_1855_),
    .D(_2060_),
    .Y(_2068_));
 OR5x2_ASAP7_75t_R _5013_ (.A(_0788_),
    .B(_1857_),
    .C(_1863_),
    .D(_2067_),
    .E(_2068_),
    .Y(_2069_));
 TAPCELL_ASAP7_75t_R PHY_121 ();
 AND4x2_ASAP7_75t_R _5015_ (.A(_1963_),
    .B(_2057_),
    .C(_2065_),
    .D(_2069_),
    .Y(_2071_));
 NAND2x2_ASAP7_75t_R _5016_ (.A(_2055_),
    .B(_2071_),
    .Y(_2072_));
 OR2x2_ASAP7_75t_R _5017_ (.A(_2053_),
    .B(_2072_),
    .Y(_2073_));
 NAND2x2_ASAP7_75t_R _5018_ (.A(net180),
    .B(_2073_),
    .Y(_3260_));
 CKINVDCx5p33_ASAP7_75t_R _5019_ (.A(_3260_),
    .Y(_3254_));
 INVx2_ASAP7_75t_R _5020_ (.A(_0179_),
    .Y(_2074_));
 AND2x2_ASAP7_75t_R _5021_ (.A(_2074_),
    .B(_1877_),
    .Y(_2075_));
 TAPCELL_ASAP7_75t_R PHY_120 ();
 AND2x2_ASAP7_75t_R _5023_ (.A(_0797_),
    .B(net180),
    .Y(_2077_));
 XNOR2x2_ASAP7_75t_R _5024_ (.A(_2075_),
    .B(_2077_),
    .Y(_3613_));
 TAPCELL_ASAP7_75t_R PHY_119 ();
 TAPCELL_ASAP7_75t_R PHY_118 ();
 TAPCELL_ASAP7_75t_R PHY_117 ();
 AND2x2_ASAP7_75t_R _5028_ (.A(_0208_),
    .B(net180),
    .Y(_2081_));
 AO21x2_ASAP7_75t_R _5029_ (.A1(net162),
    .A2(_3614_),
    .B(_2081_),
    .Y(_3616_));
 INVx3_ASAP7_75t_R _5030_ (.A(_2053_),
    .Y(_3619_));
 NAND2x2_ASAP7_75t_R _5031_ (.A(_2065_),
    .B(_2069_),
    .Y(_2082_));
 AND2x2_ASAP7_75t_R _5032_ (.A(_0211_),
    .B(net180),
    .Y(_2083_));
 XNOR2x2_ASAP7_75t_R _5033_ (.A(_2082_),
    .B(_2083_),
    .Y(_3617_));
 AND2x2_ASAP7_75t_R _5034_ (.A(_0213_),
    .B(net180),
    .Y(_2084_));
 AO21x2_ASAP7_75t_R _5035_ (.A1(net162),
    .A2(_2055_),
    .B(_2084_),
    .Y(_3283_));
 TAPCELL_ASAP7_75t_R PHY_116 ();
 OR2x2_ASAP7_75t_R _5037_ (.A(_2007_),
    .B(net222),
    .Y(_2086_));
 AND2x2_ASAP7_75t_R _5038_ (.A(_0800_),
    .B(net180),
    .Y(_2087_));
 XNOR2x2_ASAP7_75t_R _5039_ (.A(_2017_),
    .B(_2087_),
    .Y(_2088_));
 XNOR2x2_ASAP7_75t_R _5040_ (.A(_2086_),
    .B(_2088_),
    .Y(_3620_));
 AND3x2_ASAP7_75t_R _5041_ (.A(_0606_),
    .B(_1956_),
    .C(_1961_),
    .Y(_2089_));
 AO21x2_ASAP7_75t_R _5042_ (.A1(net228),
    .A2(_3236_),
    .B(_2089_),
    .Y(_3621_));
 AND2x2_ASAP7_75t_R _5043_ (.A(_0217_),
    .B(net180),
    .Y(_2090_));
 AO21x2_ASAP7_75t_R _5044_ (.A1(net162),
    .A2(_3621_),
    .B(_2090_),
    .Y(_3623_));
 INVx2_ASAP7_75t_R _5045_ (.A(_2039_),
    .Y(_3630_));
 NAND2x2_ASAP7_75t_R _5046_ (.A(_2042_),
    .B(_2046_),
    .Y(_2091_));
 AND2x2_ASAP7_75t_R _5047_ (.A(_3630_),
    .B(_2091_),
    .Y(_3626_));
 AND2x2_ASAP7_75t_R _5048_ (.A(_0802_),
    .B(net180),
    .Y(_2092_));
 AND3x2_ASAP7_75t_R _5049_ (.A(_1956_),
    .B(_1961_),
    .C(_2049_),
    .Y(_2093_));
 AO21x2_ASAP7_75t_R _5050_ (.A1(net222),
    .A2(_1972_),
    .B(_2093_),
    .Y(_2094_));
 XOR2x2_ASAP7_75t_R _5051_ (.A(_2092_),
    .B(_2094_),
    .Y(_3624_));
 OR2x2_ASAP7_75t_R _5052_ (.A(_1877_),
    .B(_1975_),
    .Y(_2095_));
 OA21x2_ASAP7_75t_R _5053_ (.A1(_2048_),
    .A2(net222),
    .B(_2095_),
    .Y(_3625_));
 AND2x2_ASAP7_75t_R _5054_ (.A(_0221_),
    .B(net180),
    .Y(_2096_));
 AO21x2_ASAP7_75t_R _5055_ (.A1(net162),
    .A2(_3625_),
    .B(_2096_),
    .Y(_3627_));
 AND2x2_ASAP7_75t_R _5056_ (.A(_0804_),
    .B(net180),
    .Y(_2097_));
 NOR2x2_ASAP7_75t_R _5057_ (.A(_1877_),
    .B(_1980_),
    .Y(_2098_));
 AO21x2_ASAP7_75t_R _5058_ (.A1(_1877_),
    .A2(_2044_),
    .B(_2098_),
    .Y(_2099_));
 XOR2x2_ASAP7_75t_R _5059_ (.A(_2097_),
    .B(_2099_),
    .Y(_3628_));
 OR2x2_ASAP7_75t_R _5060_ (.A(_2043_),
    .B(net236),
    .Y(_2100_));
 OA21x2_ASAP7_75t_R _5061_ (.A1(_1877_),
    .A2(_1935_),
    .B(_2100_),
    .Y(_3629_));
 AND2x2_ASAP7_75t_R _5062_ (.A(net162),
    .B(_3629_),
    .Y(_2101_));
 AND2x2_ASAP7_75t_R _5063_ (.A(_0225_),
    .B(net180),
    .Y(_2102_));
 OR2x2_ASAP7_75t_R _5064_ (.A(_2101_),
    .B(_2102_),
    .Y(_3631_));
 INVx2_ASAP7_75t_R _5065_ (.A(_0186_),
    .Y(_2103_));
 OR2x2_ASAP7_75t_R _5066_ (.A(_2103_),
    .B(_1864_),
    .Y(_2104_));
 OA21x2_ASAP7_75t_R _5067_ (.A1(_1877_),
    .A2(_3247_),
    .B(_2104_),
    .Y(_3637_));
 AO32x2_ASAP7_75t_R _5068_ (.A1(_1677_),
    .A2(_2056_),
    .A3(_1992_),
    .B1(_1991_),
    .B2(_1863_),
    .Y(_2105_));
 NAND2x2_ASAP7_75t_R _5069_ (.A(_2025_),
    .B(_2027_),
    .Y(_2106_));
 NOR2x2_ASAP7_75t_R _5070_ (.A(_0187_),
    .B(_2033_),
    .Y(_2107_));
 XOR2x2_ASAP7_75t_R _5071_ (.A(_0608_),
    .B(_0786_),
    .Y(_2108_));
 AND3x2_ASAP7_75t_R _5072_ (.A(_3642_),
    .B(_2107_),
    .C(_2108_),
    .Y(_2109_));
 AO22x2_ASAP7_75t_R _5073_ (.A1(_2105_),
    .A2(_2106_),
    .B1(_2109_),
    .B2(_1877_),
    .Y(_2110_));
 AND2x2_ASAP7_75t_R _5074_ (.A(_3637_),
    .B(_2110_),
    .Y(_3634_));
 AND2x2_ASAP7_75t_R _5075_ (.A(_0806_),
    .B(net180),
    .Y(_2111_));
 INVx2_ASAP7_75t_R _5076_ (.A(_2036_),
    .Y(_2112_));
 NOR2x2_ASAP7_75t_R _5077_ (.A(_1877_),
    .B(_1986_),
    .Y(_2113_));
 AO21x2_ASAP7_75t_R _5078_ (.A1(_1877_),
    .A2(_2112_),
    .B(_2113_),
    .Y(_2114_));
 XOR2x2_ASAP7_75t_R _5079_ (.A(_2111_),
    .B(_2114_),
    .Y(_3632_));
 INVx2_ASAP7_75t_R _5080_ (.A(_3245_),
    .Y(_2115_));
 INVx2_ASAP7_75t_R _5081_ (.A(_0185_),
    .Y(_2116_));
 AND2x2_ASAP7_75t_R _5082_ (.A(_2116_),
    .B(_1877_),
    .Y(_2117_));
 AO21x2_ASAP7_75t_R _5083_ (.A1(net222),
    .A2(_2115_),
    .B(_2117_),
    .Y(_3633_));
 AND2x2_ASAP7_75t_R _5084_ (.A(net162),
    .B(_3633_),
    .Y(_2118_));
 AND2x2_ASAP7_75t_R _5085_ (.A(_0229_),
    .B(net180),
    .Y(_2119_));
 OR2x2_ASAP7_75t_R _5086_ (.A(_2118_),
    .B(_2119_),
    .Y(_3635_));
 AND2x2_ASAP7_75t_R _5087_ (.A(_0808_),
    .B(net180),
    .Y(_2120_));
 OA21x2_ASAP7_75t_R _5088_ (.A1(net228),
    .A2(_2034_),
    .B(_2020_),
    .Y(_2121_));
 XNOR2x2_ASAP7_75t_R _5089_ (.A(_2120_),
    .B(_2121_),
    .Y(_3636_));
 AND2x2_ASAP7_75t_R _5090_ (.A(net162),
    .B(_3637_),
    .Y(_2122_));
 AND2x2_ASAP7_75t_R _5091_ (.A(_0233_),
    .B(net180),
    .Y(_2123_));
 OR2x2_ASAP7_75t_R _5092_ (.A(_2122_),
    .B(_2123_),
    .Y(_3639_));
 AND2x2_ASAP7_75t_R _5093_ (.A(_0810_),
    .B(net180),
    .Y(_2124_));
 OR2x2_ASAP7_75t_R _5094_ (.A(_2021_),
    .B(_2023_),
    .Y(_2125_));
 TAPCELL_ASAP7_75t_R PHY_115 ();
 OR2x2_ASAP7_75t_R _5096_ (.A(_1677_),
    .B(_2125_),
    .Y(_2126_));
 OA21x2_ASAP7_75t_R _5097_ (.A1(net221),
    .A2(_2026_),
    .B(_2126_),
    .Y(_3607_));
 AND2x2_ASAP7_75t_R _5098_ (.A(_1877_),
    .B(_2033_),
    .Y(_2127_));
 AO21x2_ASAP7_75t_R _5099_ (.A1(net228),
    .A2(_3607_),
    .B(_2127_),
    .Y(_2128_));
 XNOR2x2_ASAP7_75t_R _5100_ (.A(_2124_),
    .B(_2128_),
    .Y(_3640_));
 INVx2_ASAP7_75t_R _5101_ (.A(_0187_),
    .Y(_2129_));
 OR2x2_ASAP7_75t_R _5102_ (.A(_2129_),
    .B(net236),
    .Y(_2130_));
 OA21x2_ASAP7_75t_R _5103_ (.A1(_1877_),
    .A2(_3249_),
    .B(_2130_),
    .Y(_3641_));
 AND2x2_ASAP7_75t_R _5104_ (.A(net162),
    .B(_3641_),
    .Y(_2131_));
 AND2x2_ASAP7_75t_R _5105_ (.A(_0237_),
    .B(net180),
    .Y(_2132_));
 OR2x2_ASAP7_75t_R _5106_ (.A(_2131_),
    .B(_2132_),
    .Y(_3643_));
 INVx2_ASAP7_75t_R _5107_ (.A(_3647_),
    .Y(_3270_));
 OA21x2_ASAP7_75t_R _5108_ (.A1(_0239_),
    .A2(_3270_),
    .B(_0238_),
    .Y(_2133_));
 OA21x2_ASAP7_75t_R _5109_ (.A1(_0809_),
    .A2(_2133_),
    .B(_0236_),
    .Y(_3274_));
 OR2x2_ASAP7_75t_R _5110_ (.A(_0235_),
    .B(_0807_),
    .Y(_2134_));
 OA21x2_ASAP7_75t_R _5111_ (.A1(_0234_),
    .A2(_0807_),
    .B(_0232_),
    .Y(_2135_));
 OA21x2_ASAP7_75t_R _5112_ (.A1(_3274_),
    .A2(_2134_),
    .B(_2135_),
    .Y(_3276_));
 OA21x2_ASAP7_75t_R _5113_ (.A1(_0231_),
    .A2(_3276_),
    .B(_0230_),
    .Y(_2136_));
 OA21x2_ASAP7_75t_R _5114_ (.A1(_0805_),
    .A2(_2136_),
    .B(_0228_),
    .Y(_2137_));
 TAPCELL_ASAP7_75t_R PHY_114 ();
 OR2x2_ASAP7_75t_R _5116_ (.A(_0223_),
    .B(_0803_),
    .Y(_2138_));
 OA21x2_ASAP7_75t_R _5117_ (.A1(_0226_),
    .A2(_0803_),
    .B(_0224_),
    .Y(_2139_));
 OA21x2_ASAP7_75t_R _5118_ (.A1(_0223_),
    .A2(_2139_),
    .B(_0222_),
    .Y(_2140_));
 AND3x2_ASAP7_75t_R _5119_ (.A(_0218_),
    .B(_0220_),
    .C(_2140_),
    .Y(_2141_));
 OA31x2_ASAP7_75t_R _5120_ (.A1(_0227_),
    .A2(_2137_),
    .A3(_2138_),
    .B1(_2141_),
    .Y(_2142_));
 AO21x2_ASAP7_75t_R _5121_ (.A1(_0220_),
    .A2(_0801_),
    .B(_0219_),
    .Y(_2143_));
 AND2x2_ASAP7_75t_R _5122_ (.A(_0218_),
    .B(_2143_),
    .Y(_2144_));
 OR3x2_ASAP7_75t_R _5123_ (.A(_0215_),
    .B(_0799_),
    .C(_0798_),
    .Y(_2145_));
 OR2x2_ASAP7_75t_R _5124_ (.A(_0215_),
    .B(_0216_),
    .Y(_2146_));
 AO21x2_ASAP7_75t_R _5125_ (.A1(_0214_),
    .A2(_2146_),
    .B(_0798_),
    .Y(_2147_));
 OA31x2_ASAP7_75t_R _5126_ (.A1(_2142_),
    .A2(_2144_),
    .A3(_2145_),
    .B1(_2147_),
    .Y(_2148_));
 AND2x2_ASAP7_75t_R _5127_ (.A(_0212_),
    .B(_2148_),
    .Y(_3267_));
 AND3x2_ASAP7_75t_R _5128_ (.A(_0209_),
    .B(_0207_),
    .C(_0212_),
    .Y(_2149_));
 AND3x2_ASAP7_75t_R _5129_ (.A(_0209_),
    .B(_0207_),
    .C(_0210_),
    .Y(_2150_));
 AO21x2_ASAP7_75t_R _5130_ (.A1(_0207_),
    .A2(_0796_),
    .B(_2150_),
    .Y(_2151_));
 OR2x2_ASAP7_75t_R _5131_ (.A(_0206_),
    .B(_0795_),
    .Y(_2152_));
 AO211x2_ASAP7_75t_R _5132_ (.A1(_2148_),
    .A2(_2149_),
    .B(_2151_),
    .C(_2152_),
    .Y(_2153_));
 OA21x2_ASAP7_75t_R _5133_ (.A1(_0205_),
    .A2(_0795_),
    .B(_0204_),
    .Y(_2154_));
 AO21x2_ASAP7_75t_R _5134_ (.A1(_2153_),
    .A2(_2154_),
    .B(_0203_),
    .Y(_2155_));
 AND3x2_ASAP7_75t_R _5135_ (.A(_0199_),
    .B(_0202_),
    .C(_0794_),
    .Y(_2156_));
 AND3x2_ASAP7_75t_R _5136_ (.A(_0199_),
    .B(_0201_),
    .C(_0794_),
    .Y(_2157_));
 AO221x2_ASAP7_75t_R _5137_ (.A1(_0199_),
    .A2(_0200_),
    .B1(_2155_),
    .B2(_2156_),
    .C(_2157_),
    .Y(_2158_));
 OA21x2_ASAP7_75t_R _5138_ (.A1(_0793_),
    .A2(_2158_),
    .B(_0198_),
    .Y(_3259_));
 OR2x2_ASAP7_75t_R _5139_ (.A(_0195_),
    .B(_0197_),
    .Y(_2159_));
 OR2x2_ASAP7_75t_R _5140_ (.A(_0793_),
    .B(_2159_),
    .Y(_2160_));
 OA222x2_ASAP7_75t_R _5141_ (.A1(_0196_),
    .A2(_0195_),
    .B1(_0198_),
    .B2(_2159_),
    .C1(_2160_),
    .C2(_2158_),
    .Y(_2161_));
 AND3x2_ASAP7_75t_R _5142_ (.A(_0193_),
    .B(_0792_),
    .C(_0791_),
    .Y(_2162_));
 AND3x2_ASAP7_75t_R _5143_ (.A(_0193_),
    .B(_0194_),
    .C(_0791_),
    .Y(_2163_));
 AO221x2_ASAP7_75t_R _5144_ (.A1(_0192_),
    .A2(_0791_),
    .B1(_2161_),
    .B2(_2162_),
    .C(_2163_),
    .Y(_3256_));
 OA21x2_ASAP7_75t_R _5145_ (.A1(_0191_),
    .A2(_3256_),
    .B(_0190_),
    .Y(_2164_));
 OA21x2_ASAP7_75t_R _5146_ (.A1(_0189_),
    .A2(_2164_),
    .B(_0790_),
    .Y(_3255_));
 AND2x2_ASAP7_75t_R _5147_ (.A(_0792_),
    .B(_2161_),
    .Y(_3257_));
 AND2x2_ASAP7_75t_R _5148_ (.A(_2153_),
    .B(_2154_),
    .Y(_3263_));
 OR3x2_ASAP7_75t_R _5149_ (.A(_0227_),
    .B(_2137_),
    .C(_2138_),
    .Y(_2165_));
 AO21x2_ASAP7_75t_R _5150_ (.A1(_2165_),
    .A2(_2140_),
    .B(_0801_),
    .Y(_2166_));
 AND2x2_ASAP7_75t_R _5151_ (.A(_0220_),
    .B(_2166_),
    .Y(_3282_));
 OA21x2_ASAP7_75t_R _5152_ (.A1(_0227_),
    .A2(_2137_),
    .B(_0226_),
    .Y(_2167_));
 OA21x2_ASAP7_75t_R _5153_ (.A1(_0803_),
    .A2(_2167_),
    .B(_0224_),
    .Y(_3280_));
 TAPCELL_ASAP7_75t_R PHY_113 ();
 INVx2_ASAP7_75t_R _5155_ (.A(_0259_),
    .Y(\__st_2[6] ));
 INVx2_ASAP7_75t_R _5156_ (.A(_0563_),
    .Y(\__st_2[4] ));
 TAPCELL_ASAP7_75t_R PHY_112 ();
 OA21x2_ASAP7_75t_R _5158_ (.A1(_0258_),
    .A2(_3293_),
    .B(_0257_),
    .Y(_2170_));
 OA21x2_ASAP7_75t_R _5159_ (.A1(_0816_),
    .A2(_2170_),
    .B(_0256_),
    .Y(_2171_));
 OR3x2_ASAP7_75t_R _5160_ (.A(_0562_),
    .B(_0563_),
    .C(_2171_),
    .Y(_2172_));
 OR3x2_ASAP7_75t_R _5161_ (.A(_0255_),
    .B(_0259_),
    .C(_2172_),
    .Y(_2173_));
 AO21x2_ASAP7_75t_R _5162_ (.A1(_0254_),
    .A2(_2173_),
    .B(_0253_),
    .Y(_2174_));
 AO21x2_ASAP7_75t_R _5163_ (.A1(_0252_),
    .A2(_2174_),
    .B(_0251_),
    .Y(_2175_));
 AND2x2_ASAP7_75t_R _5164_ (.A(_0250_),
    .B(_2175_),
    .Y(_3290_));
 OA21x2_ASAP7_75t_R _5165_ (.A1(_0249_),
    .A2(_3290_),
    .B(_0248_),
    .Y(_2176_));
 OA21x2_ASAP7_75t_R _5166_ (.A1(_0815_),
    .A2(_2176_),
    .B(_0247_),
    .Y(_3288_));
 OA21x2_ASAP7_75t_R _5167_ (.A1(_0246_),
    .A2(_3288_),
    .B(_0245_),
    .Y(_2177_));
 OA21x2_ASAP7_75t_R _5168_ (.A1(_0814_),
    .A2(_2177_),
    .B(_0244_),
    .Y(_3286_));
 INVx2_ASAP7_75t_R _5169_ (.A(_2172_),
    .Y(_3648_));
 INVx2_ASAP7_75t_R _5170_ (.A(_0557_),
    .Y(\__st_2[13] ));
 INVx2_ASAP7_75t_R _5171_ (.A(_3287_),
    .Y(\__st_2[12] ));
 INVx2_ASAP7_75t_R _5172_ (.A(_0558_),
    .Y(\__st_2[11] ));
 INVx2_ASAP7_75t_R _5173_ (.A(_3289_),
    .Y(\__st_2[10] ));
 INVx2_ASAP7_75t_R _5174_ (.A(_0559_),
    .Y(\__st_2[9] ));
 INVx2_ASAP7_75t_R _5175_ (.A(_0560_),
    .Y(\__st_2[8] ));
 INVx2_ASAP7_75t_R _5176_ (.A(_0561_),
    .Y(\__st_2[7] ));
 INVx2_ASAP7_75t_R _5177_ (.A(_0564_),
    .Y(\__st_2[3] ));
 INVx2_ASAP7_75t_R _5178_ (.A(_3292_),
    .Y(\__st_2[2] ));
 INVx2_ASAP7_75t_R _5179_ (.A(_0565_),
    .Y(\__st_2[1] ));
 INVx2_ASAP7_75t_R _5180_ (.A(_0566_),
    .Y(\__st_2[0] ));
 INVx3_ASAP7_75t_R _5181_ (.A(_0822_),
    .Y(_3655_));
 AND4x2_ASAP7_75t_R _5182_ (.A(_3289_),
    .B(_0559_),
    .C(_0560_),
    .D(_0561_),
    .Y(_2178_));
 AND4x2_ASAP7_75t_R _5183_ (.A(_3285_),
    .B(_0557_),
    .C(_3287_),
    .D(_0558_),
    .Y(_2179_));
 OA21x2_ASAP7_75t_R _5184_ (.A1(_0259_),
    .A2(_0562_),
    .B(_0564_),
    .Y(_2180_));
 AND3x2_ASAP7_75t_R _5185_ (.A(_2178_),
    .B(_2179_),
    .C(_2180_),
    .Y(_2181_));
 OA21x2_ASAP7_75t_R _5186_ (.A1(_0563_),
    .A2(_0564_),
    .B(_0562_),
    .Y(_2182_));
 OA211x2_ASAP7_75t_R _5187_ (.A1(_0259_),
    .A2(_2182_),
    .B(_2179_),
    .C(_2178_),
    .Y(_2183_));
 TAPCELL_ASAP7_75t_R PHY_111 ();
 INVx2_ASAP7_75t_R _5189_ (.A(_2183_),
    .Y(_2185_));
 OR2x2_ASAP7_75t_R _5190_ (.A(_3292_),
    .B(_2185_),
    .Y(_3654_));
 AND2x2_ASAP7_75t_R _5191_ (.A(_3655_),
    .B(_3654_),
    .Y(_2186_));
 NOR2x2_ASAP7_75t_R _5192_ (.A(_2181_),
    .B(_2186_),
    .Y(_3653_));
 AND2x6_ASAP7_75t_R _5193_ (.A(_2178_),
    .B(_2179_),
    .Y(_2187_));
 OA21x2_ASAP7_75t_R _5194_ (.A1(_0259_),
    .A2(_0562_),
    .B(_0563_),
    .Y(_2188_));
 NAND2x2_ASAP7_75t_R _5195_ (.A(_2187_),
    .B(_2188_),
    .Y(_3652_));
 INVx2_ASAP7_75t_R _5196_ (.A(_0562_),
    .Y(_2189_));
 AND4x2_ASAP7_75t_R _5197_ (.A(_0259_),
    .B(_2189_),
    .C(_2178_),
    .D(_2179_),
    .Y(_2190_));
 AO21x2_ASAP7_75t_R _5198_ (.A1(_3653_),
    .A2(_3652_),
    .B(_2190_),
    .Y(_3651_));
 TAPCELL_ASAP7_75t_R PHY_110 ();
 INVx2_ASAP7_75t_R _5200_ (.A(_0821_),
    .Y(_2192_));
 XNOR2x2_ASAP7_75t_R _5201_ (.A(_2192_),
    .B(_2181_),
    .Y(_2193_));
 OR2x6_ASAP7_75t_R _5202_ (.A(_0820_),
    .B(_2193_),
    .Y(_2194_));
 TAPCELL_ASAP7_75t_R PHY_109 ();
 XNOR2x2_ASAP7_75t_R _5204_ (.A(_0819_),
    .B(_2190_),
    .Y(_2196_));
 TAPCELL_ASAP7_75t_R PHY_108 ();
 NOR2x2_ASAP7_75t_R _5206_ (.A(_3655_),
    .B(_2183_),
    .Y(_2198_));
 TAPCELL_ASAP7_75t_R PHY_107 ();
 INVx2_ASAP7_75t_R _5208_ (.A(_0818_),
    .Y(_2200_));
 OR2x2_ASAP7_75t_R _5209_ (.A(_0265_),
    .B(_2200_),
    .Y(_2201_));
 OR4x2_ASAP7_75t_R _5210_ (.A(_2194_),
    .B(_2196_),
    .C(_2198_),
    .D(_2201_),
    .Y(_2202_));
 TAPCELL_ASAP7_75t_R PHY_106 ();
 INVx3_ASAP7_75t_R _5212_ (.A(_2202_),
    .Y(_3337_));
 TAPCELL_ASAP7_75t_R PHY_105 ();
 TAPCELL_ASAP7_75t_R PHY_104 ();
 TAPCELL_ASAP7_75t_R PHY_103 ();
 TAPCELL_ASAP7_75t_R PHY_102 ();
 OA21x2_ASAP7_75t_R _5217_ (.A1(_0259_),
    .A2(_2182_),
    .B(\__st_2[0] ),
    .Y(_2207_));
 AND2x6_ASAP7_75t_R _5218_ (.A(_2187_),
    .B(_2207_),
    .Y(_2208_));
 CKINVDCx16_ASAP7_75t_R _5219_ (.A(_2208_),
    .Y(_2209_));
 TAPCELL_ASAP7_75t_R PHY_101 ();
 TAPCELL_ASAP7_75t_R PHY_100 ();
 TAPCELL_ASAP7_75t_R PHY_99 ();
 OA21x2_ASAP7_75t_R _5223_ (.A1(net48),
    .A2(_2209_),
    .B(_2193_),
    .Y(_2213_));
 INVx11_ASAP7_75t_R _5224_ (.A(net40),
    .Y(_2214_));
 OA21x2_ASAP7_75t_R _5225_ (.A1(_3655_),
    .A2(_2183_),
    .B(_2214_),
    .Y(_2215_));
 XOR2x2_ASAP7_75t_R _5226_ (.A(_0819_),
    .B(_2190_),
    .Y(_2216_));
 INVx2_ASAP7_75t_R _5227_ (.A(_0265_),
    .Y(_2217_));
 AND2x2_ASAP7_75t_R _5228_ (.A(_2217_),
    .B(_0818_),
    .Y(_2218_));
 AND2x2_ASAP7_75t_R _5229_ (.A(_2216_),
    .B(_2218_),
    .Y(_2219_));
 OA211x2_ASAP7_75t_R _5230_ (.A1(net45),
    .A2(_2213_),
    .B(_2215_),
    .C(_2219_),
    .Y(_2220_));
 TAPCELL_ASAP7_75t_R PHY_98 ();
 CKINVDCx12_ASAP7_75t_R _5232_ (.A(net44),
    .Y(_2221_));
 CKINVDCx10_ASAP7_75t_R _5233_ (.A(net49),
    .Y(_2222_));
 AND2x2_ASAP7_75t_R _5234_ (.A(_2221_),
    .B(_2222_),
    .Y(_2223_));
 TAPCELL_ASAP7_75t_R PHY_97 ();
 AND2x4_ASAP7_75t_R _5236_ (.A(_2193_),
    .B(_2208_),
    .Y(_2225_));
 AND2x2_ASAP7_75t_R _5237_ (.A(_2223_),
    .B(_2225_),
    .Y(_2226_));
 AND2x2_ASAP7_75t_R _5238_ (.A(_2193_),
    .B(_2209_),
    .Y(_2227_));
 OA21x2_ASAP7_75t_R _5239_ (.A1(net48),
    .A2(_2227_),
    .B(net45),
    .Y(_2228_));
 TAPCELL_ASAP7_75t_R PHY_96 ();
 OA21x2_ASAP7_75t_R _5241_ (.A1(_2226_),
    .A2(_2228_),
    .B(_2214_),
    .Y(_2230_));
 XNOR2x2_ASAP7_75t_R _5242_ (.A(_0821_),
    .B(_2181_),
    .Y(_2231_));
 TAPCELL_ASAP7_75t_R PHY_95 ();
 TAPCELL_ASAP7_75t_R PHY_94 ();
 OR2x2_ASAP7_75t_R _5245_ (.A(net40),
    .B(_2209_),
    .Y(_2234_));
 AND2x2_ASAP7_75t_R _5246_ (.A(_0266_),
    .B(net40),
    .Y(_2235_));
 AO21x2_ASAP7_75t_R _5247_ (.A1(net48),
    .A2(_2234_),
    .B(_2235_),
    .Y(_2236_));
 AND2x2_ASAP7_75t_R _5248_ (.A(_2231_),
    .B(_2236_),
    .Y(_2237_));
 OR2x6_ASAP7_75t_R _5249_ (.A(_3655_),
    .B(_2183_),
    .Y(_2238_));
 AND2x2_ASAP7_75t_R _5250_ (.A(_2238_),
    .B(_2218_),
    .Y(_2239_));
 OA211x2_ASAP7_75t_R _5251_ (.A1(_2230_),
    .A2(_2237_),
    .B(_2216_),
    .C(_2239_),
    .Y(_2240_));
 TAPCELL_ASAP7_75t_R PHY_93 ();
 TAPCELL_ASAP7_75t_R PHY_92 ();
 TAPCELL_ASAP7_75t_R PHY_91 ();
 OR2x2_ASAP7_75t_R _5255_ (.A(net48),
    .B(_2193_),
    .Y(_2243_));
 AND2x2_ASAP7_75t_R _5256_ (.A(_2222_),
    .B(_2231_),
    .Y(_2244_));
 AND2x2_ASAP7_75t_R _5257_ (.A(net48),
    .B(_2193_),
    .Y(_2245_));
 OR3x2_ASAP7_75t_R _5258_ (.A(_0266_),
    .B(_2244_),
    .C(_2245_),
    .Y(_2246_));
 OA211x2_ASAP7_75t_R _5259_ (.A1(_2221_),
    .A2(_2243_),
    .B(_2246_),
    .C(_2238_),
    .Y(_2247_));
 TAPCELL_ASAP7_75t_R PHY_90 ();
 AND2x2_ASAP7_75t_R _5261_ (.A(_2221_),
    .B(net49),
    .Y(_2249_));
 AND2x6_ASAP7_75t_R _5262_ (.A(_2231_),
    .B(_2208_),
    .Y(_2250_));
 TAPCELL_ASAP7_75t_R PHY_89 ();
 OR2x4_ASAP7_75t_R _5264_ (.A(_2231_),
    .B(_2208_),
    .Y(_2252_));
 OR2x2_ASAP7_75t_R _5265_ (.A(_2193_),
    .B(_2209_),
    .Y(_2253_));
 OA211x2_ASAP7_75t_R _5266_ (.A1(net48),
    .A2(_2252_),
    .B(_2253_),
    .C(_2238_),
    .Y(_2254_));
 TAPCELL_ASAP7_75t_R PHY_88 ();
 OA21x2_ASAP7_75t_R _5268_ (.A1(_0266_),
    .A2(_2193_),
    .B(_2209_),
    .Y(_2256_));
 OR2x2_ASAP7_75t_R _5269_ (.A(_2222_),
    .B(_2256_),
    .Y(_2257_));
 TAPCELL_ASAP7_75t_R PHY_87 ();
 TAPCELL_ASAP7_75t_R PHY_86 ();
 AO221x2_ASAP7_75t_R _5272_ (.A1(_2249_),
    .A2(_2250_),
    .B1(_2254_),
    .B2(_2257_),
    .C(net40),
    .Y(_2260_));
 OA211x2_ASAP7_75t_R _5273_ (.A1(_2214_),
    .A2(_2247_),
    .B(_2260_),
    .C(_2219_),
    .Y(_2261_));
 TAPCELL_ASAP7_75t_R PHY_85 ();
 OR2x2_ASAP7_75t_R _5275_ (.A(_2221_),
    .B(_2231_),
    .Y(_2262_));
 AND2x2_ASAP7_75t_R _5276_ (.A(_2222_),
    .B(net40),
    .Y(_2263_));
 OA21x2_ASAP7_75t_R _5277_ (.A1(_2216_),
    .A2(_2209_),
    .B(_2214_),
    .Y(_2264_));
 AO33x2_ASAP7_75t_R _5278_ (.A1(_2216_),
    .A2(_2262_),
    .A3(_2263_),
    .B1(_2264_),
    .B2(_2243_),
    .B3(_2252_),
    .Y(_2265_));
 AND2x2_ASAP7_75t_R _5279_ (.A(_2214_),
    .B(_2231_),
    .Y(_2266_));
 AND2x2_ASAP7_75t_R _5280_ (.A(_2266_),
    .B(_2196_),
    .Y(_2267_));
 AND2x2_ASAP7_75t_R _5281_ (.A(net48),
    .B(_0820_),
    .Y(_2268_));
 AND3x2_ASAP7_75t_R _5282_ (.A(_2216_),
    .B(_2227_),
    .C(_2268_),
    .Y(_2269_));
 OA21x2_ASAP7_75t_R _5283_ (.A1(_2267_),
    .A2(_2269_),
    .B(net45),
    .Y(_2270_));
 OA21x2_ASAP7_75t_R _5284_ (.A1(_2265_),
    .A2(_2270_),
    .B(_2239_),
    .Y(_2271_));
 TAPCELL_ASAP7_75t_R PHY_84 ();
 AO21x2_ASAP7_75t_R _5286_ (.A1(_0820_),
    .A2(_2208_),
    .B(_2215_),
    .Y(_2272_));
 AND2x2_ASAP7_75t_R _5287_ (.A(net45),
    .B(net48),
    .Y(_2273_));
 AND2x2_ASAP7_75t_R _5288_ (.A(_2193_),
    .B(_2273_),
    .Y(_2274_));
 AO21x2_ASAP7_75t_R _5289_ (.A1(_2272_),
    .A2(_2274_),
    .B(_2196_),
    .Y(_2275_));
 OA21x2_ASAP7_75t_R _5290_ (.A1(_2214_),
    .A2(_2209_),
    .B(_2231_),
    .Y(_2276_));
 NOR2x2_ASAP7_75t_R _5291_ (.A(_2192_),
    .B(_2180_),
    .Y(_2277_));
 AND2x2_ASAP7_75t_R _5292_ (.A(_2192_),
    .B(_2180_),
    .Y(_2278_));
 OA211x2_ASAP7_75t_R _5293_ (.A1(_2277_),
    .A2(_2278_),
    .B(_2187_),
    .C(_2207_),
    .Y(_2279_));
 OR3x2_ASAP7_75t_R _5294_ (.A(_0267_),
    .B(_0820_),
    .C(_2279_),
    .Y(_2280_));
 OA21x2_ASAP7_75t_R _5295_ (.A1(_2221_),
    .A2(_2209_),
    .B(_2238_),
    .Y(_2281_));
 OA211x2_ASAP7_75t_R _5296_ (.A1(_2222_),
    .A2(_2276_),
    .B(_2280_),
    .C(_2281_),
    .Y(_2282_));
 OA21x2_ASAP7_75t_R _5297_ (.A1(_3655_),
    .A2(_2183_),
    .B(_2222_),
    .Y(_2283_));
 OA21x2_ASAP7_75t_R _5298_ (.A1(_2208_),
    .A2(_2283_),
    .B(_2221_),
    .Y(_2284_));
 AND3x2_ASAP7_75t_R _5299_ (.A(_2238_),
    .B(_2209_),
    .C(_2273_),
    .Y(_2285_));
 OR4x2_ASAP7_75t_R _5300_ (.A(_2193_),
    .B(_2216_),
    .C(_2284_),
    .D(_2285_),
    .Y(_2286_));
 OA21x2_ASAP7_75t_R _5301_ (.A1(_3655_),
    .A2(_2183_),
    .B(net45),
    .Y(_2287_));
 OA21x2_ASAP7_75t_R _5302_ (.A1(_2231_),
    .A2(_2287_),
    .B(_2214_),
    .Y(_2288_));
 OA21x2_ASAP7_75t_R _5303_ (.A1(_2216_),
    .A2(_2288_),
    .B(_2218_),
    .Y(_2289_));
 OA211x2_ASAP7_75t_R _5304_ (.A1(_2275_),
    .A2(_2282_),
    .B(_2286_),
    .C(_2289_),
    .Y(_2290_));
 TAPCELL_ASAP7_75t_R PHY_83 ();
 AND3x2_ASAP7_75t_R _5306_ (.A(net49),
    .B(_2187_),
    .C(_2207_),
    .Y(_2291_));
 AO21x2_ASAP7_75t_R _5307_ (.A1(_2209_),
    .A2(_2283_),
    .B(_2291_),
    .Y(_2292_));
 AND2x2_ASAP7_75t_R _5308_ (.A(_2231_),
    .B(_2292_),
    .Y(_2293_));
 AND2x2_ASAP7_75t_R _5309_ (.A(_2193_),
    .B(_2238_),
    .Y(_2294_));
 OA21x2_ASAP7_75t_R _5310_ (.A1(_2250_),
    .A2(_2294_),
    .B(_2221_),
    .Y(_2295_));
 OA21x2_ASAP7_75t_R _5311_ (.A1(_2293_),
    .A2(_2295_),
    .B(_2214_),
    .Y(_2296_));
 TAPCELL_ASAP7_75t_R PHY_82 ();
 OR2x2_ASAP7_75t_R _5313_ (.A(net48),
    .B(_2209_),
    .Y(_2298_));
 AND3x2_ASAP7_75t_R _5314_ (.A(_2231_),
    .B(_2238_),
    .C(_2298_),
    .Y(_2299_));
 TAPCELL_ASAP7_75t_R PHY_81 ();
 AO21x2_ASAP7_75t_R _5316_ (.A1(_2235_),
    .A2(_2299_),
    .B(_2216_),
    .Y(_2301_));
 OR2x2_ASAP7_75t_R _5317_ (.A(_2214_),
    .B(_2231_),
    .Y(_2302_));
 AND3x2_ASAP7_75t_R _5318_ (.A(_0266_),
    .B(_2234_),
    .C(_2302_),
    .Y(_2303_));
 OR2x2_ASAP7_75t_R _5319_ (.A(net48),
    .B(_0820_),
    .Y(_2304_));
 OR2x2_ASAP7_75t_R _5320_ (.A(_2193_),
    .B(_2208_),
    .Y(_2305_));
 OR2x2_ASAP7_75t_R _5321_ (.A(_2222_),
    .B(_2231_),
    .Y(_2306_));
 OA211x2_ASAP7_75t_R _5322_ (.A1(_2304_),
    .A2(_2305_),
    .B(_2221_),
    .C(_2306_),
    .Y(_2307_));
 OR2x2_ASAP7_75t_R _5323_ (.A(net49),
    .B(_2214_),
    .Y(_2308_));
 AO21x2_ASAP7_75t_R _5324_ (.A1(_2231_),
    .A2(_2308_),
    .B(_2209_),
    .Y(_2309_));
 OA211x2_ASAP7_75t_R _5325_ (.A1(_2303_),
    .A2(_2307_),
    .B(_2239_),
    .C(_2309_),
    .Y(_2310_));
 AND2x2_ASAP7_75t_R _5326_ (.A(net49),
    .B(_2214_),
    .Y(_2311_));
 AO21x2_ASAP7_75t_R _5327_ (.A1(_2221_),
    .A2(_2311_),
    .B(_2235_),
    .Y(_2312_));
 AO21x2_ASAP7_75t_R _5328_ (.A1(_2225_),
    .A2(_2312_),
    .B(_2196_),
    .Y(_2313_));
 AND2x2_ASAP7_75t_R _5329_ (.A(_2218_),
    .B(_2313_),
    .Y(_2314_));
 OA22x2_ASAP7_75t_R _5330_ (.A1(_2296_),
    .A2(_2301_),
    .B1(_2310_),
    .B2(_2314_),
    .Y(_2315_));
 TAPCELL_ASAP7_75t_R PHY_80 ();
 TAPCELL_ASAP7_75t_R PHY_79 ();
 AND2x2_ASAP7_75t_R _5333_ (.A(net40),
    .B(_2231_),
    .Y(_2317_));
 AO21x2_ASAP7_75t_R _5334_ (.A1(_2214_),
    .A2(_2231_),
    .B(net48),
    .Y(_2318_));
 AO221x2_ASAP7_75t_R _5335_ (.A1(_2223_),
    .A2(_2317_),
    .B1(_2318_),
    .B2(_0266_),
    .C(_2245_),
    .Y(_2319_));
 AND2x2_ASAP7_75t_R _5336_ (.A(_2221_),
    .B(_2214_),
    .Y(_2320_));
 AO21x2_ASAP7_75t_R _5337_ (.A1(_2305_),
    .A2(_2320_),
    .B(_2225_),
    .Y(_2321_));
 AND2x2_ASAP7_75t_R _5338_ (.A(_2222_),
    .B(_2208_),
    .Y(_2322_));
 OA21x2_ASAP7_75t_R _5339_ (.A1(_2193_),
    .A2(_2322_),
    .B(_2235_),
    .Y(_2323_));
 AO221x2_ASAP7_75t_R _5340_ (.A1(_2209_),
    .A2(_2319_),
    .B1(_2321_),
    .B2(_2222_),
    .C(_2323_),
    .Y(_2324_));
 AO21x2_ASAP7_75t_R _5341_ (.A1(_2194_),
    .A2(_2302_),
    .B(_0266_),
    .Y(_2325_));
 OR2x2_ASAP7_75t_R _5342_ (.A(net49),
    .B(_2231_),
    .Y(_2326_));
 OA21x2_ASAP7_75t_R _5343_ (.A1(_2221_),
    .A2(net40),
    .B(_2209_),
    .Y(_2327_));
 OR2x2_ASAP7_75t_R _5344_ (.A(_2221_),
    .B(_2193_),
    .Y(_2328_));
 OA22x2_ASAP7_75t_R _5345_ (.A1(_2326_),
    .A2(_2327_),
    .B1(_2328_),
    .B2(_2322_),
    .Y(_2329_));
 TAPCELL_ASAP7_75t_R PHY_78 ();
 OA211x2_ASAP7_75t_R _5347_ (.A1(_0266_),
    .A2(net48),
    .B(_2218_),
    .C(_2208_),
    .Y(_2331_));
 AO32x2_ASAP7_75t_R _5348_ (.A1(_2239_),
    .A2(_2325_),
    .A3(_2329_),
    .B1(_2331_),
    .B2(_2266_),
    .Y(_2332_));
 AO32x2_ASAP7_75t_R _5349_ (.A1(_2238_),
    .A2(_2219_),
    .A3(_2324_),
    .B1(_2332_),
    .B2(_2196_),
    .Y(_2333_));
 TAPCELL_ASAP7_75t_R PHY_77 ();
 OR2x2_ASAP7_75t_R _5351_ (.A(_2221_),
    .B(_2222_),
    .Y(_2334_));
 OR4x2_ASAP7_75t_R _5352_ (.A(_2200_),
    .B(_2196_),
    .C(_2198_),
    .D(_2334_),
    .Y(_2335_));
 OA21x2_ASAP7_75t_R _5353_ (.A1(_2194_),
    .A2(_2335_),
    .B(_2201_),
    .Y(_2336_));
 OA21x2_ASAP7_75t_R _5354_ (.A1(net40),
    .A2(_2209_),
    .B(_2221_),
    .Y(_2337_));
 AO21x2_ASAP7_75t_R _5355_ (.A1(_2187_),
    .A2(_2207_),
    .B(_0820_),
    .Y(_2338_));
 OA211x2_ASAP7_75t_R _5356_ (.A1(_2209_),
    .A2(_2308_),
    .B(_2338_),
    .C(net44),
    .Y(_2339_));
 AO21x2_ASAP7_75t_R _5357_ (.A1(_2302_),
    .A2(_2337_),
    .B(_2339_),
    .Y(_2340_));
 AO221x2_ASAP7_75t_R _5358_ (.A1(_0822_),
    .A2(_2185_),
    .B1(_2305_),
    .B2(_0266_),
    .C(_2222_),
    .Y(_2341_));
 OA211x2_ASAP7_75t_R _5359_ (.A1(_2198_),
    .A2(_2340_),
    .B(_2341_),
    .C(_2194_),
    .Y(_2342_));
 INVx2_ASAP7_75t_R _5360_ (.A(_2292_),
    .Y(_2343_));
 OA21x2_ASAP7_75t_R _5361_ (.A1(net45),
    .A2(_2343_),
    .B(_2266_),
    .Y(_2344_));
 OR4x2_ASAP7_75t_R _5362_ (.A(_2216_),
    .B(_2336_),
    .C(_2342_),
    .D(_2344_),
    .Y(_2345_));
 AND2x2_ASAP7_75t_R _5363_ (.A(_2193_),
    .B(_2311_),
    .Y(_2346_));
 OR3x2_ASAP7_75t_R _5364_ (.A(_2221_),
    .B(_2263_),
    .C(_2346_),
    .Y(_2347_));
 OA211x2_ASAP7_75t_R _5365_ (.A1(_0266_),
    .A2(_2317_),
    .B(_2347_),
    .C(_2209_),
    .Y(_2348_));
 OA211x2_ASAP7_75t_R _5366_ (.A1(_2253_),
    .A2(_2304_),
    .B(_2216_),
    .C(_2238_),
    .Y(_2349_));
 OR2x2_ASAP7_75t_R _5367_ (.A(net44),
    .B(_2231_),
    .Y(_2350_));
 AO21x2_ASAP7_75t_R _5368_ (.A1(_2209_),
    .A2(_2304_),
    .B(_2350_),
    .Y(_2351_));
 NAND2x2_ASAP7_75t_R _5369_ (.A(_2349_),
    .B(_2351_),
    .Y(_2352_));
 OA21x2_ASAP7_75t_R _5370_ (.A1(_2348_),
    .A2(_2352_),
    .B(_2217_),
    .Y(_2353_));
 OR2x2_ASAP7_75t_R _5371_ (.A(_2336_),
    .B(_2353_),
    .Y(_2354_));
 NAND2x2_ASAP7_75t_R _5372_ (.A(_2345_),
    .B(_2354_),
    .Y(_3348_));
 AO21x2_ASAP7_75t_R _5373_ (.A1(_2231_),
    .A2(_2208_),
    .B(_2222_),
    .Y(_2355_));
 AO21x2_ASAP7_75t_R _5374_ (.A1(_2243_),
    .A2(_2355_),
    .B(_2198_),
    .Y(_2356_));
 OR2x2_ASAP7_75t_R _5375_ (.A(_2221_),
    .B(_2209_),
    .Y(_2357_));
 OA21x2_ASAP7_75t_R _5376_ (.A1(net48),
    .A2(_2198_),
    .B(_2193_),
    .Y(_2358_));
 OA21x2_ASAP7_75t_R _5377_ (.A1(_2357_),
    .A2(_2358_),
    .B(_0820_),
    .Y(_2359_));
 OA21x2_ASAP7_75t_R _5378_ (.A1(net45),
    .A2(_2356_),
    .B(_2359_),
    .Y(_2360_));
 OR2x2_ASAP7_75t_R _5379_ (.A(_2222_),
    .B(_2208_),
    .Y(_2361_));
 OA21x2_ASAP7_75t_R _5380_ (.A1(net44),
    .A2(_2361_),
    .B(_2298_),
    .Y(_2362_));
 AND2x2_ASAP7_75t_R _5381_ (.A(_2214_),
    .B(_2193_),
    .Y(_2363_));
 OA21x2_ASAP7_75t_R _5382_ (.A1(_2198_),
    .A2(_2362_),
    .B(_2363_),
    .Y(_2364_));
 OR2x2_ASAP7_75t_R _5383_ (.A(_2198_),
    .B(_2208_),
    .Y(_2365_));
 OA21x2_ASAP7_75t_R _5384_ (.A1(net45),
    .A2(_2365_),
    .B(_2266_),
    .Y(_2366_));
 OR4x2_ASAP7_75t_R _5385_ (.A(_2216_),
    .B(_2360_),
    .C(_2364_),
    .D(_2366_),
    .Y(_2367_));
 AND2x2_ASAP7_75t_R _5386_ (.A(_2231_),
    .B(_2209_),
    .Y(_2368_));
 OA211x2_ASAP7_75t_R _5387_ (.A1(_2368_),
    .A2(_2363_),
    .B(net45),
    .C(_2222_),
    .Y(_2369_));
 AND3x2_ASAP7_75t_R _5388_ (.A(_2221_),
    .B(_0820_),
    .C(_2193_),
    .Y(_2370_));
 OA211x2_ASAP7_75t_R _5389_ (.A1(_2266_),
    .A2(_2370_),
    .B(_2209_),
    .C(_2222_),
    .Y(_2371_));
 AO21x2_ASAP7_75t_R _5390_ (.A1(net40),
    .A2(_2250_),
    .B(_2346_),
    .Y(_2372_));
 AND2x2_ASAP7_75t_R _5391_ (.A(_2221_),
    .B(_2372_),
    .Y(_2373_));
 AND2x2_ASAP7_75t_R _5392_ (.A(_2252_),
    .B(_2268_),
    .Y(_2374_));
 AND2x2_ASAP7_75t_R _5393_ (.A(net45),
    .B(_2225_),
    .Y(_2375_));
 OR4x2_ASAP7_75t_R _5394_ (.A(_2196_),
    .B(_2198_),
    .C(_2374_),
    .D(_2375_),
    .Y(_2376_));
 OR4x2_ASAP7_75t_R _5395_ (.A(_2369_),
    .B(_2371_),
    .C(_2373_),
    .D(_2376_),
    .Y(_2377_));
 AND2x2_ASAP7_75t_R _5396_ (.A(_2252_),
    .B(_2273_),
    .Y(_2378_));
 INVx2_ASAP7_75t_R _5397_ (.A(_2378_),
    .Y(_2379_));
 AND2x2_ASAP7_75t_R _5398_ (.A(_0818_),
    .B(_2216_),
    .Y(_2380_));
 OA211x2_ASAP7_75t_R _5399_ (.A1(_2231_),
    .A2(_2273_),
    .B(_2380_),
    .C(_2215_),
    .Y(_2381_));
 NAND2x2_ASAP7_75t_R _5400_ (.A(_2379_),
    .B(_2381_),
    .Y(_2382_));
 AO32x2_ASAP7_75t_R _5401_ (.A1(_2217_),
    .A2(_2367_),
    .A3(_2377_),
    .B1(_2201_),
    .B2(_2382_),
    .Y(_2383_));
 TAPCELL_ASAP7_75t_R PHY_76 ();
 INVx4_ASAP7_75t_R _5403_ (.A(_2383_),
    .Y(_3325_));
 TAPCELL_ASAP7_75t_R PHY_75 ();
 TAPCELL_ASAP7_75t_R PHY_74 ();
 TAPCELL_ASAP7_75t_R PHY_73 ();
 AO21x2_ASAP7_75t_R _5407_ (.A1(net49),
    .A2(_2209_),
    .B(_2193_),
    .Y(_2386_));
 TAPCELL_ASAP7_75t_R PHY_72 ();
 TAPCELL_ASAP7_75t_R PHY_71 ();
 AND2x2_ASAP7_75t_R _5410_ (.A(_0266_),
    .B(_2222_),
    .Y(_2389_));
 AO21x2_ASAP7_75t_R _5411_ (.A1(_2221_),
    .A2(_2386_),
    .B(_2389_),
    .Y(_2390_));
 AO21x2_ASAP7_75t_R _5412_ (.A1(_2238_),
    .A2(_2390_),
    .B(_2279_),
    .Y(_2391_));
 TAPCELL_ASAP7_75t_R PHY_70 ();
 TAPCELL_ASAP7_75t_R PHY_69 ();
 AO21x2_ASAP7_75t_R _5415_ (.A1(_2231_),
    .A2(_2285_),
    .B(_2214_),
    .Y(_2394_));
 OA211x2_ASAP7_75t_R _5416_ (.A1(_0820_),
    .A2(_2391_),
    .B(_2394_),
    .C(_2380_),
    .Y(_2395_));
 AO21x2_ASAP7_75t_R _5417_ (.A1(_2209_),
    .A2(_2328_),
    .B(net49),
    .Y(_2396_));
 OR2x2_ASAP7_75t_R _5418_ (.A(_0266_),
    .B(_2222_),
    .Y(_2397_));
 AND2x2_ASAP7_75t_R _5419_ (.A(_2238_),
    .B(_2397_),
    .Y(_2398_));
 AO221x2_ASAP7_75t_R _5420_ (.A1(_2225_),
    .A2(_2249_),
    .B1(_2396_),
    .B2(_2398_),
    .C(_2214_),
    .Y(_2399_));
 AND2x2_ASAP7_75t_R _5421_ (.A(_2221_),
    .B(_2208_),
    .Y(_2400_));
 AO21x2_ASAP7_75t_R _5422_ (.A1(net49),
    .A2(_2209_),
    .B(_2400_),
    .Y(_2401_));
 AO21x2_ASAP7_75t_R _5423_ (.A1(_2238_),
    .A2(_2401_),
    .B(_2194_),
    .Y(_2402_));
 MAJx2_ASAP7_75t_R _5424_ (.A(net44),
    .B(_2222_),
    .C(_2209_),
    .Y(_2403_));
 AO32x2_ASAP7_75t_R _5425_ (.A1(_2187_),
    .A2(_2207_),
    .A3(_2249_),
    .B1(_2403_),
    .B2(_2238_),
    .Y(_2404_));
 OR3x2_ASAP7_75t_R _5426_ (.A(_0820_),
    .B(_2231_),
    .C(_2404_),
    .Y(_2405_));
 AND3x2_ASAP7_75t_R _5427_ (.A(_2399_),
    .B(_2402_),
    .C(_2405_),
    .Y(_2406_));
 OA21x2_ASAP7_75t_R _5428_ (.A1(_2231_),
    .A2(_2322_),
    .B(net44),
    .Y(_2407_));
 AND3x2_ASAP7_75t_R _5429_ (.A(_2221_),
    .B(_2222_),
    .C(_2209_),
    .Y(_2408_));
 OA21x2_ASAP7_75t_R _5430_ (.A1(_2407_),
    .A2(_2408_),
    .B(_2238_),
    .Y(_2409_));
 AO21x2_ASAP7_75t_R _5431_ (.A1(_2249_),
    .A2(_2250_),
    .B(_2409_),
    .Y(_2410_));
 MAJx2_ASAP7_75t_R _5432_ (.A(net49),
    .B(_2209_),
    .C(_2363_),
    .Y(_2411_));
 AND2x2_ASAP7_75t_R _5433_ (.A(_2214_),
    .B(_2208_),
    .Y(_2412_));
 OA211x2_ASAP7_75t_R _5434_ (.A1(_2193_),
    .A2(_2412_),
    .B(_2221_),
    .C(_2222_),
    .Y(_2413_));
 AO21x2_ASAP7_75t_R _5435_ (.A1(net44),
    .A2(_2411_),
    .B(_2413_),
    .Y(_2414_));
 AO221x2_ASAP7_75t_R _5436_ (.A1(net40),
    .A2(_2410_),
    .B1(_2414_),
    .B2(_2238_),
    .C(_2216_),
    .Y(_2415_));
 OA21x2_ASAP7_75t_R _5437_ (.A1(_2196_),
    .A2(_2406_),
    .B(_2415_),
    .Y(_2416_));
 OA22x2_ASAP7_75t_R _5438_ (.A1(_2218_),
    .A2(_2395_),
    .B1(_2416_),
    .B2(_0265_),
    .Y(_2417_));
 TAPCELL_ASAP7_75t_R PHY_68 ();
 INVx2_ASAP7_75t_R _5440_ (.A(_2417_),
    .Y(_3310_));
 AO21x2_ASAP7_75t_R _5441_ (.A1(net45),
    .A2(_2243_),
    .B(_2346_),
    .Y(_2418_));
 OR2x2_ASAP7_75t_R _5442_ (.A(_2214_),
    .B(_2250_),
    .Y(_2419_));
 AO21x2_ASAP7_75t_R _5443_ (.A1(net40),
    .A2(_2252_),
    .B(net45),
    .Y(_2420_));
 OA211x2_ASAP7_75t_R _5444_ (.A1(_2221_),
    .A2(_2419_),
    .B(_2420_),
    .C(_2222_),
    .Y(_2421_));
 AO221x2_ASAP7_75t_R _5445_ (.A1(net45),
    .A2(_2363_),
    .B1(_2418_),
    .B2(_2209_),
    .C(_2421_),
    .Y(_2422_));
 AO32x2_ASAP7_75t_R _5446_ (.A1(_2221_),
    .A2(_2250_),
    .A3(_2304_),
    .B1(_2422_),
    .B2(_2238_),
    .Y(_2423_));
 AO32x2_ASAP7_75t_R _5447_ (.A1(_0820_),
    .A2(_2193_),
    .A3(_2273_),
    .B1(_2250_),
    .B2(_2222_),
    .Y(_2424_));
 AO21x2_ASAP7_75t_R _5448_ (.A1(_2252_),
    .A2(_2243_),
    .B(net45),
    .Y(_2425_));
 INVx2_ASAP7_75t_R _5449_ (.A(_2425_),
    .Y(_2426_));
 OA211x2_ASAP7_75t_R _5450_ (.A1(_2424_),
    .A2(_2426_),
    .B(_2196_),
    .C(_2238_),
    .Y(_2427_));
 AO21x2_ASAP7_75t_R _5451_ (.A1(_2216_),
    .A2(_2423_),
    .B(_2427_),
    .Y(_2428_));
 AO21x2_ASAP7_75t_R _5452_ (.A1(_2238_),
    .A2(_2334_),
    .B(_2208_),
    .Y(_2429_));
 AO21x2_ASAP7_75t_R _5453_ (.A1(_2231_),
    .A2(_2429_),
    .B(_2214_),
    .Y(_2430_));
 AND2x2_ASAP7_75t_R _5454_ (.A(_2216_),
    .B(_2430_),
    .Y(_2431_));
 AO21x2_ASAP7_75t_R _5455_ (.A1(net45),
    .A2(_2252_),
    .B(_2222_),
    .Y(_2432_));
 OA211x2_ASAP7_75t_R _5456_ (.A1(net45),
    .A2(_2368_),
    .B(_2253_),
    .C(_2238_),
    .Y(_2433_));
 AO221x2_ASAP7_75t_R _5457_ (.A1(_2249_),
    .A2(_2250_),
    .B1(_2432_),
    .B2(_2433_),
    .C(_0820_),
    .Y(_2434_));
 AO21x2_ASAP7_75t_R _5458_ (.A1(_2431_),
    .A2(_2434_),
    .B(_2217_),
    .Y(_2435_));
 OA211x2_ASAP7_75t_R _5459_ (.A1(_0265_),
    .A2(_2428_),
    .B(_2435_),
    .C(_0818_),
    .Y(_2436_));
 TAPCELL_ASAP7_75t_R PHY_67 ();
 INVx2_ASAP7_75t_R _5461_ (.A(_2436_),
    .Y(_3328_));
 TAPCELL_ASAP7_75t_R PHY_66 ();
 OA22x2_ASAP7_75t_R _5463_ (.A1(_2208_),
    .A2(_2308_),
    .B1(_2311_),
    .B2(net44),
    .Y(_2438_));
 AO21x2_ASAP7_75t_R _5464_ (.A1(_2234_),
    .A2(_2438_),
    .B(_2231_),
    .Y(_2439_));
 AO21x2_ASAP7_75t_R _5465_ (.A1(_2222_),
    .A2(_2338_),
    .B(_2328_),
    .Y(_2440_));
 OA211x2_ASAP7_75t_R _5466_ (.A1(_2209_),
    .A2(_2397_),
    .B(_2196_),
    .C(_2238_),
    .Y(_2441_));
 OA21x2_ASAP7_75t_R _5467_ (.A1(_2194_),
    .A2(_2404_),
    .B(_2216_),
    .Y(_2442_));
 TAPCELL_ASAP7_75t_R PHY_65 ();
 OA21x2_ASAP7_75t_R _5469_ (.A1(net48),
    .A2(_2208_),
    .B(_2231_),
    .Y(_2444_));
 AO21x2_ASAP7_75t_R _5470_ (.A1(_2209_),
    .A2(_2235_),
    .B(_2444_),
    .Y(_2445_));
 INVx2_ASAP7_75t_R _5471_ (.A(_2445_),
    .Y(_2446_));
 OR2x2_ASAP7_75t_R _5472_ (.A(net48),
    .B(_2198_),
    .Y(_2447_));
 OA21x2_ASAP7_75t_R _5473_ (.A1(_2252_),
    .A2(_2447_),
    .B(_2234_),
    .Y(_2448_));
 OA222x2_ASAP7_75t_R _5474_ (.A1(_0820_),
    .A2(_2213_),
    .B1(_2446_),
    .B2(_2198_),
    .C1(_2448_),
    .C2(_0266_),
    .Y(_2449_));
 INVx2_ASAP7_75t_R _5475_ (.A(_2449_),
    .Y(_2450_));
 AO32x2_ASAP7_75t_R _5476_ (.A1(_2439_),
    .A2(_2440_),
    .A3(_2441_),
    .B1(_2442_),
    .B2(_2450_),
    .Y(_2451_));
 AO221x2_ASAP7_75t_R _5477_ (.A1(_2209_),
    .A2(_2283_),
    .B1(_2279_),
    .B2(net48),
    .C(_2221_),
    .Y(_2452_));
 AO221x2_ASAP7_75t_R _5478_ (.A1(_2231_),
    .A2(_2208_),
    .B1(_2294_),
    .B2(net48),
    .C(_0266_),
    .Y(_2453_));
 AO21x2_ASAP7_75t_R _5479_ (.A1(net48),
    .A2(_2227_),
    .B(_2250_),
    .Y(_2454_));
 AND2x2_ASAP7_75t_R _5480_ (.A(net40),
    .B(_2454_),
    .Y(_2455_));
 OR2x2_ASAP7_75t_R _5481_ (.A(_2244_),
    .B(_2455_),
    .Y(_2456_));
 AO32x2_ASAP7_75t_R _5482_ (.A1(_2214_),
    .A2(_2452_),
    .A3(_2453_),
    .B1(_2287_),
    .B2(_2456_),
    .Y(_2457_));
 AO21x2_ASAP7_75t_R _5483_ (.A1(_2216_),
    .A2(_2457_),
    .B(_2217_),
    .Y(_2458_));
 OA211x2_ASAP7_75t_R _5484_ (.A1(_0265_),
    .A2(_2451_),
    .B(_2458_),
    .C(_0818_),
    .Y(_2459_));
 TAPCELL_ASAP7_75t_R PHY_64 ();
 AO21x2_ASAP7_75t_R _5486_ (.A1(_2238_),
    .A2(_2227_),
    .B(_2250_),
    .Y(_2460_));
 AO21x2_ASAP7_75t_R _5487_ (.A1(_2231_),
    .A2(_2238_),
    .B(net45),
    .Y(_2461_));
 OA211x2_ASAP7_75t_R _5488_ (.A1(_2221_),
    .A2(_2460_),
    .B(_2461_),
    .C(net48),
    .Y(_2462_));
 NOR2x2_ASAP7_75t_R _5489_ (.A(_2214_),
    .B(_2462_),
    .Y(_2463_));
 OR3x2_ASAP7_75t_R _5490_ (.A(_2198_),
    .B(_2389_),
    .C(_2400_),
    .Y(_2464_));
 OA21x2_ASAP7_75t_R _5491_ (.A1(_2397_),
    .A2(_2365_),
    .B(_2357_),
    .Y(_2465_));
 INVx2_ASAP7_75t_R _5492_ (.A(_2380_),
    .Y(_2466_));
 AO221x2_ASAP7_75t_R _5493_ (.A1(_2363_),
    .A2(_2464_),
    .B1(_2465_),
    .B2(_2266_),
    .C(_2466_),
    .Y(_2467_));
 OA21x2_ASAP7_75t_R _5494_ (.A1(_2463_),
    .A2(_2467_),
    .B(_2201_),
    .Y(_2468_));
 INVx2_ASAP7_75t_R _5495_ (.A(_2389_),
    .Y(_2469_));
 AO21x2_ASAP7_75t_R _5496_ (.A1(_2194_),
    .A2(_2208_),
    .B(_2469_),
    .Y(_2470_));
 OR2x2_ASAP7_75t_R _5497_ (.A(_2221_),
    .B(_2326_),
    .Y(_2471_));
 OA21x2_ASAP7_75t_R _5498_ (.A1(net44),
    .A2(_2305_),
    .B(_2471_),
    .Y(_2472_));
 OA21x2_ASAP7_75t_R _5499_ (.A1(net49),
    .A2(_2234_),
    .B(_2361_),
    .Y(_2473_));
 AND2x2_ASAP7_75t_R _5500_ (.A(_2221_),
    .B(_2194_),
    .Y(_2474_));
 OR2x2_ASAP7_75t_R _5501_ (.A(_2222_),
    .B(_2209_),
    .Y(_2475_));
 OA222x2_ASAP7_75t_R _5502_ (.A1(_2214_),
    .A2(_2472_),
    .B1(_2473_),
    .B2(_2350_),
    .C1(_2474_),
    .C2(_2475_),
    .Y(_2476_));
 AO32x2_ASAP7_75t_R _5503_ (.A1(_2196_),
    .A2(_2470_),
    .A3(_2476_),
    .B1(_2185_),
    .B2(_0822_),
    .Y(_2477_));
 OA21x2_ASAP7_75t_R _5504_ (.A1(_2263_),
    .A2(_2311_),
    .B(_2227_),
    .Y(_2478_));
 OA21x2_ASAP7_75t_R _5505_ (.A1(_2374_),
    .A2(_2478_),
    .B(net45),
    .Y(_2479_));
 OA21x2_ASAP7_75t_R _5506_ (.A1(_2225_),
    .A2(_2368_),
    .B(_2214_),
    .Y(_2480_));
 OA21x2_ASAP7_75t_R _5507_ (.A1(_2455_),
    .A2(_2480_),
    .B(_2221_),
    .Y(_2481_));
 OA21x2_ASAP7_75t_R _5508_ (.A1(_2479_),
    .A2(_2481_),
    .B(_2216_),
    .Y(_2482_));
 OA21x2_ASAP7_75t_R _5509_ (.A1(_2477_),
    .A2(_2482_),
    .B(_2217_),
    .Y(_2483_));
 OR2x2_ASAP7_75t_R _5510_ (.A(_2468_),
    .B(_2483_),
    .Y(_2484_));
 TAPCELL_ASAP7_75t_R PHY_63 ();
 INVx2_ASAP7_75t_R _5512_ (.A(_2484_),
    .Y(_3658_));
 AND2x2_ASAP7_75t_R _5513_ (.A(_2231_),
    .B(_2334_),
    .Y(_2485_));
 OA211x2_ASAP7_75t_R _5514_ (.A1(_2274_),
    .A2(_2485_),
    .B(_2238_),
    .C(_2209_),
    .Y(_2486_));
 AND3x2_ASAP7_75t_R _5515_ (.A(net45),
    .B(net48),
    .C(_2209_),
    .Y(_2487_));
 OA21x2_ASAP7_75t_R _5516_ (.A1(_2322_),
    .A2(_2487_),
    .B(_2238_),
    .Y(_2488_));
 OR3x2_ASAP7_75t_R _5517_ (.A(_2194_),
    .B(_2284_),
    .C(_2488_),
    .Y(_2489_));
 OA211x2_ASAP7_75t_R _5518_ (.A1(net45),
    .A2(_2198_),
    .B(_2357_),
    .C(_2363_),
    .Y(_2490_));
 NOR2x2_ASAP7_75t_R _5519_ (.A(_2466_),
    .B(_2490_),
    .Y(_2491_));
 OA211x2_ASAP7_75t_R _5520_ (.A1(_2214_),
    .A2(_2486_),
    .B(_2489_),
    .C(_2491_),
    .Y(_2492_));
 AO21x2_ASAP7_75t_R _5521_ (.A1(_0820_),
    .A2(_2294_),
    .B(_2250_),
    .Y(_2493_));
 OR2x2_ASAP7_75t_R _5522_ (.A(_2208_),
    .B(_2287_),
    .Y(_2494_));
 AO221x2_ASAP7_75t_R _5523_ (.A1(_2225_),
    .A2(_2320_),
    .B1(_2494_),
    .B2(_2317_),
    .C(_2216_),
    .Y(_2495_));
 AO21x2_ASAP7_75t_R _5524_ (.A1(net48),
    .A2(_2493_),
    .B(_2495_),
    .Y(_2496_));
 AO21x2_ASAP7_75t_R _5525_ (.A1(net49),
    .A2(_2231_),
    .B(net44),
    .Y(_2497_));
 OR3x2_ASAP7_75t_R _5526_ (.A(_2221_),
    .B(_2193_),
    .C(_2311_),
    .Y(_2498_));
 AO21x2_ASAP7_75t_R _5527_ (.A1(net44),
    .A2(_2214_),
    .B(_2193_),
    .Y(_2499_));
 AO32x2_ASAP7_75t_R _5528_ (.A1(_2209_),
    .A2(_2497_),
    .A3(_2498_),
    .B1(_2499_),
    .B2(_2322_),
    .Y(_2500_));
 AO221x2_ASAP7_75t_R _5529_ (.A1(_2193_),
    .A2(_2412_),
    .B1(_2500_),
    .B2(_2238_),
    .C(_2196_),
    .Y(_2501_));
 AO21x2_ASAP7_75t_R _5530_ (.A1(_2496_),
    .A2(_2501_),
    .B(_0265_),
    .Y(_2502_));
 OA21x2_ASAP7_75t_R _5531_ (.A1(_2218_),
    .A2(_2492_),
    .B(_2502_),
    .Y(_3669_));
 INVx2_ASAP7_75t_R _5532_ (.A(_3667_),
    .Y(_3309_));
 OA21x2_ASAP7_75t_R _5533_ (.A1(_0282_),
    .A2(_3309_),
    .B(_0281_),
    .Y(_2503_));
 OA21x2_ASAP7_75t_R _5534_ (.A1(_0827_),
    .A2(_2503_),
    .B(_0280_),
    .Y(_2504_));
 OA21x2_ASAP7_75t_R _5535_ (.A1(_0279_),
    .A2(_2504_),
    .B(_0278_),
    .Y(_2505_));
 OA21x2_ASAP7_75t_R _5536_ (.A1(_0826_),
    .A2(_2505_),
    .B(_0277_),
    .Y(_3303_));
 OA21x2_ASAP7_75t_R _5537_ (.A1(_0276_),
    .A2(_3303_),
    .B(_0275_),
    .Y(_2506_));
 OA21x2_ASAP7_75t_R _5538_ (.A1(_0825_),
    .A2(_2506_),
    .B(_0274_),
    .Y(_3300_));
 OA21x2_ASAP7_75t_R _5539_ (.A1(_0273_),
    .A2(_3300_),
    .B(_0272_),
    .Y(_2507_));
 OA21x2_ASAP7_75t_R _5540_ (.A1(_0824_),
    .A2(_2507_),
    .B(_0271_),
    .Y(_3297_));
 OA21x2_ASAP7_75t_R _5541_ (.A1(_0270_),
    .A2(_3297_),
    .B(_0269_),
    .Y(_2508_));
 OR2x2_ASAP7_75t_R _5542_ (.A(_0823_),
    .B(_2508_),
    .Y(_2509_));
 NAND2x2_ASAP7_75t_R _5543_ (.A(_0268_),
    .B(_2509_),
    .Y(_3661_));
 AND3x2_ASAP7_75t_R _5544_ (.A(_2220_),
    .B(_2240_),
    .C(_3661_),
    .Y(_3659_));
 OR2x2_ASAP7_75t_R _5545_ (.A(_0284_),
    .B(net229),
    .Y(_2510_));
 INVx2_ASAP7_75t_R _5546_ (.A(_2510_),
    .Y(_3670_));
 INVx2_ASAP7_75t_R _5547_ (.A(_2220_),
    .Y(_3295_));
 XOR2x2_ASAP7_75t_R _5548_ (.A(_0829_),
    .B(_2220_),
    .Y(_2511_));
 NOR2x2_ASAP7_75t_R _5549_ (.A(net229),
    .B(_2511_),
    .Y(_3660_));
 OR2x4_ASAP7_75t_R _5550_ (.A(_0287_),
    .B(net229),
    .Y(_2512_));
 TAPCELL_ASAP7_75t_R PHY_62 ();
 INVx2_ASAP7_75t_R _5552_ (.A(_2512_),
    .Y(_3316_));
 INVx2_ASAP7_75t_R _5553_ (.A(_2261_),
    .Y(_3298_));
 INVx2_ASAP7_75t_R _5554_ (.A(_2271_),
    .Y(_3296_));
 INVx2_ASAP7_75t_R _5555_ (.A(_2290_),
    .Y(_3301_));
 INVx2_ASAP7_75t_R _5556_ (.A(_2315_),
    .Y(_3299_));
 INVx2_ASAP7_75t_R _5557_ (.A(_3348_),
    .Y(_3302_));
 AND2x2_ASAP7_75t_R _5558_ (.A(_0656_),
    .B(net38),
    .Y(_2513_));
 AO21x2_ASAP7_75t_R _5559_ (.A1(_1508_),
    .A2(_3325_),
    .B(_2513_),
    .Y(_3668_));
 INVx2_ASAP7_75t_R _5560_ (.A(_3668_),
    .Y(_3329_));
 AND2x2_ASAP7_75t_R _5561_ (.A(_0657_),
    .B(net38),
    .Y(_2514_));
 AO21x2_ASAP7_75t_R _5562_ (.A1(_1508_),
    .A2(_2417_),
    .B(_2514_),
    .Y(_2515_));
 INVx2_ASAP7_75t_R _5563_ (.A(_2515_),
    .Y(_3331_));
 INVx2_ASAP7_75t_R _5564_ (.A(_3677_),
    .Y(_3330_));
 OA21x2_ASAP7_75t_R _5565_ (.A1(_0305_),
    .A2(_3330_),
    .B(_0304_),
    .Y(_2516_));
 OA21x2_ASAP7_75t_R _5566_ (.A1(_0835_),
    .A2(_2516_),
    .B(_0303_),
    .Y(_2517_));
 OA21x2_ASAP7_75t_R _5567_ (.A1(_0302_),
    .A2(_2517_),
    .B(_0301_),
    .Y(_2518_));
 OA21x2_ASAP7_75t_R _5568_ (.A1(_0834_),
    .A2(_2518_),
    .B(_0299_),
    .Y(_2519_));
 OA21x2_ASAP7_75t_R _5569_ (.A1(_0297_),
    .A2(_2519_),
    .B(_0296_),
    .Y(_2520_));
 OR3x2_ASAP7_75t_R _5570_ (.A(_0294_),
    .B(_0833_),
    .C(_0832_),
    .Y(_2521_));
 OR3x2_ASAP7_75t_R _5571_ (.A(_0294_),
    .B(_0295_),
    .C(_0832_),
    .Y(_2522_));
 OA211x2_ASAP7_75t_R _5572_ (.A1(_0293_),
    .A2(_0832_),
    .B(_2522_),
    .C(_0292_),
    .Y(_2523_));
 OA21x2_ASAP7_75t_R _5573_ (.A1(_2520_),
    .A2(_2521_),
    .B(_2523_),
    .Y(_2524_));
 OR2x2_ASAP7_75t_R _5574_ (.A(_0291_),
    .B(_0831_),
    .Y(_2525_));
 OA21x2_ASAP7_75t_R _5575_ (.A1(_0290_),
    .A2(_0831_),
    .B(_0830_),
    .Y(_2526_));
 OA21x2_ASAP7_75t_R _5576_ (.A1(_2524_),
    .A2(_2525_),
    .B(_2526_),
    .Y(_3314_));
 INVx2_ASAP7_75t_R _5577_ (.A(_0659_),
    .Y(_2527_));
 OR3x2_ASAP7_75t_R _5578_ (.A(_2527_),
    .B(_1598_),
    .C(_1674_),
    .Y(_2528_));
 OA21x2_ASAP7_75t_R _5579_ (.A1(_1677_),
    .A2(_2512_),
    .B(_2528_),
    .Y(_2529_));
 TAPCELL_ASAP7_75t_R PHY_61 ();
 INVx2_ASAP7_75t_R _5581_ (.A(_0661_),
    .Y(_2530_));
 AND2x2_ASAP7_75t_R _5582_ (.A(net221),
    .B(_3329_),
    .Y(_2531_));
 AO21x2_ASAP7_75t_R _5583_ (.A1(_2530_),
    .A2(_1677_),
    .B(_2531_),
    .Y(_2532_));
 TAPCELL_ASAP7_75t_R PHY_60 ();
 OA21x2_ASAP7_75t_R _5585_ (.A1(_0331_),
    .A2(_3352_),
    .B(_0330_),
    .Y(_2533_));
 OA21x2_ASAP7_75t_R _5586_ (.A1(_0842_),
    .A2(_2533_),
    .B(_0329_),
    .Y(_2534_));
 OA21x2_ASAP7_75t_R _5587_ (.A1(_0328_),
    .A2(_2534_),
    .B(_0327_),
    .Y(_2535_));
 OA21x2_ASAP7_75t_R _5588_ (.A1(_0841_),
    .A2(_2535_),
    .B(_0325_),
    .Y(_2536_));
 OA21x2_ASAP7_75t_R _5589_ (.A1(_0323_),
    .A2(_2536_),
    .B(_0322_),
    .Y(_2537_));
 OA21x2_ASAP7_75t_R _5590_ (.A1(_0840_),
    .A2(_2537_),
    .B(_0320_),
    .Y(_2538_));
 OA21x2_ASAP7_75t_R _5591_ (.A1(_0318_),
    .A2(_2538_),
    .B(_0317_),
    .Y(_2539_));
 OA21x2_ASAP7_75t_R _5592_ (.A1(_0839_),
    .A2(_2539_),
    .B(_0315_),
    .Y(_2540_));
 OA21x2_ASAP7_75t_R _5593_ (.A1(_0313_),
    .A2(_2540_),
    .B(_0312_),
    .Y(_2541_));
 OA21x2_ASAP7_75t_R _5594_ (.A1(_0838_),
    .A2(_2541_),
    .B(_0837_),
    .Y(_3336_));
 AO21x2_ASAP7_75t_R _5595_ (.A1(_1927_),
    .A2(_1855_),
    .B(_2510_),
    .Y(_2542_));
 OA21x2_ASAP7_75t_R _5596_ (.A1(_0307_),
    .A2(net219),
    .B(_2542_),
    .Y(_2543_));
 INVx2_ASAP7_75t_R _5597_ (.A(_2543_),
    .Y(_3680_));
 INVx2_ASAP7_75t_R _5598_ (.A(_2529_),
    .Y(_3338_));
 INVx2_ASAP7_75t_R _5599_ (.A(_0311_),
    .Y(_2544_));
 AND2x2_ASAP7_75t_R _5600_ (.A(net229),
    .B(_2220_),
    .Y(_2545_));
 AO21x2_ASAP7_75t_R _5601_ (.A1(_0650_),
    .A2(net223),
    .B(_2545_),
    .Y(_3318_));
 OR2x2_ASAP7_75t_R _5602_ (.A(_1677_),
    .B(_3318_),
    .Y(_2546_));
 OA21x2_ASAP7_75t_R _5603_ (.A1(_2544_),
    .A2(net219),
    .B(_2546_),
    .Y(_2547_));
 TAPCELL_ASAP7_75t_R PHY_59 ();
 NAND2x2_ASAP7_75t_R _5605_ (.A(net222),
    .B(_2547_),
    .Y(_2548_));
 OA21x2_ASAP7_75t_R _5606_ (.A1(_0334_),
    .A2(net222),
    .B(_2548_),
    .Y(_3692_));
 INVx2_ASAP7_75t_R _5607_ (.A(_0316_),
    .Y(_2549_));
 AND2x2_ASAP7_75t_R _5608_ (.A(_0652_),
    .B(net223),
    .Y(_2550_));
 AO21x2_ASAP7_75t_R _5609_ (.A1(net229),
    .A2(_2261_),
    .B(_2550_),
    .Y(_2551_));
 TAPCELL_ASAP7_75t_R PHY_58 ();
 OR2x2_ASAP7_75t_R _5611_ (.A(_1677_),
    .B(_2551_),
    .Y(_2552_));
 OA21x2_ASAP7_75t_R _5612_ (.A1(_2549_),
    .A2(net219),
    .B(_2552_),
    .Y(_2553_));
 TAPCELL_ASAP7_75t_R PHY_57 ();
 NAND2x2_ASAP7_75t_R _5614_ (.A(net222),
    .B(_2553_),
    .Y(_2554_));
 OA21x2_ASAP7_75t_R _5615_ (.A1(_0336_),
    .A2(net222),
    .B(_2554_),
    .Y(_3696_));
 INVx2_ASAP7_75t_R _5616_ (.A(_0321_),
    .Y(_2555_));
 OR2x2_ASAP7_75t_R _5617_ (.A(_2555_),
    .B(net219),
    .Y(_2556_));
 AND2x2_ASAP7_75t_R _5618_ (.A(net229),
    .B(_2290_),
    .Y(_2557_));
 AO21x2_ASAP7_75t_R _5619_ (.A1(_0654_),
    .A2(net223),
    .B(_2557_),
    .Y(_2558_));
 TAPCELL_ASAP7_75t_R PHY_56 ();
 OR2x2_ASAP7_75t_R _5621_ (.A(_1677_),
    .B(_2558_),
    .Y(_2559_));
 NAND2x2_ASAP7_75t_R _5622_ (.A(_2556_),
    .B(_2559_),
    .Y(_2560_));
 OR2x2_ASAP7_75t_R _5623_ (.A(_0338_),
    .B(net222),
    .Y(_2561_));
 OA21x2_ASAP7_75t_R _5624_ (.A1(_1877_),
    .A2(_2560_),
    .B(_2561_),
    .Y(_3700_));
 INVx2_ASAP7_75t_R _5625_ (.A(_0326_),
    .Y(_2562_));
 INVx2_ASAP7_75t_R _5626_ (.A(_0300_),
    .Y(_2563_));
 OR2x2_ASAP7_75t_R _5627_ (.A(_2563_),
    .B(_1508_),
    .Y(_2564_));
 OA21x2_ASAP7_75t_R _5628_ (.A1(net233),
    .A2(_2333_),
    .B(_2564_),
    .Y(_3326_));
 AND2x2_ASAP7_75t_R _5629_ (.A(net219),
    .B(_3326_),
    .Y(_2565_));
 AO21x2_ASAP7_75t_R _5630_ (.A1(_2562_),
    .A2(_1677_),
    .B(_2565_),
    .Y(_2566_));
 TAPCELL_ASAP7_75t_R PHY_55 ();
 NOR2x2_ASAP7_75t_R _5632_ (.A(_1877_),
    .B(_2566_),
    .Y(_2567_));
 AO21x2_ASAP7_75t_R _5633_ (.A1(_0340_),
    .A2(_1877_),
    .B(_2567_),
    .Y(_3704_));
 INVx2_ASAP7_75t_R _5634_ (.A(_0666_),
    .Y(_2568_));
 OR2x2_ASAP7_75t_R _5635_ (.A(_2568_),
    .B(net236),
    .Y(_2569_));
 OA21x2_ASAP7_75t_R _5636_ (.A1(_1877_),
    .A2(_2532_),
    .B(_2569_),
    .Y(_3708_));
 OR2x2_ASAP7_75t_R _5637_ (.A(_0662_),
    .B(net221),
    .Y(_2570_));
 OA21x2_ASAP7_75t_R _5638_ (.A1(_1677_),
    .A2(_2515_),
    .B(_2570_),
    .Y(_3354_));
 INVx2_ASAP7_75t_R _5639_ (.A(_0341_),
    .Y(_2571_));
 AND2x2_ASAP7_75t_R _5640_ (.A(_2571_),
    .B(_1877_),
    .Y(_2572_));
 AO21x2_ASAP7_75t_R _5641_ (.A1(_1864_),
    .A2(_3354_),
    .B(_2572_),
    .Y(_2573_));
 INVx2_ASAP7_75t_R _5642_ (.A(_2573_),
    .Y(_3711_));
 INVx2_ASAP7_75t_R _5643_ (.A(_0342_),
    .Y(_2574_));
 AND2x2_ASAP7_75t_R _5644_ (.A(_2574_),
    .B(_1877_),
    .Y(_2575_));
 INVx2_ASAP7_75t_R _5645_ (.A(_0332_),
    .Y(_2576_));
 INVx2_ASAP7_75t_R _5646_ (.A(_0306_),
    .Y(_2577_));
 AND2x2_ASAP7_75t_R _5647_ (.A(_2577_),
    .B(net38),
    .Y(_2578_));
 AO21x2_ASAP7_75t_R _5648_ (.A1(_1508_),
    .A2(_2436_),
    .B(_2578_),
    .Y(_3679_));
 OR2x2_ASAP7_75t_R _5649_ (.A(_1677_),
    .B(_3679_),
    .Y(_2579_));
 OA211x2_ASAP7_75t_R _5650_ (.A1(_2576_),
    .A2(net219),
    .B(_1864_),
    .C(_2579_),
    .Y(_2580_));
 NOR2x2_ASAP7_75t_R _5651_ (.A(_2575_),
    .B(_2580_),
    .Y(_3712_));
 XNOR2x2_ASAP7_75t_R _5652_ (.A(_0825_),
    .B(_0653_),
    .Y(_2581_));
 AND2x2_ASAP7_75t_R _5653_ (.A(net233),
    .B(_2581_),
    .Y(_2582_));
 AO21x2_ASAP7_75t_R _5654_ (.A1(net229),
    .A2(_2271_),
    .B(_2582_),
    .Y(_2583_));
 TAPCELL_ASAP7_75t_R PHY_54 ();
 NOR2x2_ASAP7_75t_R _5656_ (.A(_2558_),
    .B(_2583_),
    .Y(_2584_));
 XOR2x2_ASAP7_75t_R _5657_ (.A(_0319_),
    .B(_0833_),
    .Y(_2585_));
 INVx2_ASAP7_75t_R _5658_ (.A(_2585_),
    .Y(_2586_));
 AND4x2_ASAP7_75t_R _5659_ (.A(_0321_),
    .B(_1927_),
    .C(_1855_),
    .D(_2586_),
    .Y(_2587_));
 AO21x2_ASAP7_75t_R _5660_ (.A1(net219),
    .A2(_2584_),
    .B(_2587_),
    .Y(_2588_));
 XOR2x2_ASAP7_75t_R _5661_ (.A(_0324_),
    .B(_0834_),
    .Y(_2589_));
 NOR2x2_ASAP7_75t_R _5662_ (.A(_2562_),
    .B(_2589_),
    .Y(_2590_));
 XNOR2x2_ASAP7_75t_R _5663_ (.A(_0314_),
    .B(_0832_),
    .Y(_2591_));
 AND2x2_ASAP7_75t_R _5664_ (.A(_0316_),
    .B(_2591_),
    .Y(_2592_));
 XNOR2x2_ASAP7_75t_R _5665_ (.A(_0824_),
    .B(_0651_),
    .Y(_2593_));
 AND2x2_ASAP7_75t_R _5666_ (.A(net233),
    .B(_2593_),
    .Y(_2594_));
 AO21x2_ASAP7_75t_R _5667_ (.A1(net229),
    .A2(_2240_),
    .B(_2594_),
    .Y(_2595_));
 TAPCELL_ASAP7_75t_R PHY_53 ();
 NOR2x2_ASAP7_75t_R _5669_ (.A(_2551_),
    .B(_2595_),
    .Y(_2596_));
 XOR2x2_ASAP7_75t_R _5670_ (.A(_0298_),
    .B(_0826_),
    .Y(_2597_));
 INVx2_ASAP7_75t_R _5671_ (.A(_2597_),
    .Y(_2598_));
 AND3x2_ASAP7_75t_R _5672_ (.A(_0300_),
    .B(net223),
    .C(_2598_),
    .Y(_2599_));
 NOR3x2_ASAP7_75t_R _5673_ (.B(_2315_),
    .C(_2333_),
    .Y(_2600_),
    .A(net223));
 OA22x2_ASAP7_75t_R _5674_ (.A1(_1598_),
    .A2(net226),
    .B1(_2599_),
    .B2(_2600_),
    .Y(_2601_));
 AO32x2_ASAP7_75t_R _5675_ (.A1(_1677_),
    .A2(_2590_),
    .A3(_2592_),
    .B1(_2596_),
    .B2(_2601_),
    .Y(_2602_));
 XNOR2x2_ASAP7_75t_R _5676_ (.A(_0823_),
    .B(_0649_),
    .Y(_2603_));
 NOR2x2_ASAP7_75t_R _5677_ (.A(_0650_),
    .B(_2603_),
    .Y(_2604_));
 AND3x2_ASAP7_75t_R _5678_ (.A(net229),
    .B(_2202_),
    .C(_3295_),
    .Y(_2605_));
 AO21x2_ASAP7_75t_R _5679_ (.A1(net223),
    .A2(_2604_),
    .B(_2605_),
    .Y(_2606_));
 OA21x2_ASAP7_75t_R _5680_ (.A1(_1598_),
    .A2(net226),
    .B(_2606_),
    .Y(_2607_));
 XOR2x2_ASAP7_75t_R _5681_ (.A(_0310_),
    .B(_0831_),
    .Y(_2608_));
 INVx2_ASAP7_75t_R _5682_ (.A(_2608_),
    .Y(_2609_));
 AND4x2_ASAP7_75t_R _5683_ (.A(_0311_),
    .B(_1927_),
    .C(_1855_),
    .D(_2609_),
    .Y(_2610_));
 INVx2_ASAP7_75t_R _5684_ (.A(_0343_),
    .Y(_3709_));
 OA21x2_ASAP7_75t_R _5685_ (.A1(_2607_),
    .A2(_2610_),
    .B(_3709_),
    .Y(_2611_));
 XOR2x2_ASAP7_75t_R _5686_ (.A(_0827_),
    .B(_0655_),
    .Y(_2612_));
 AND2x2_ASAP7_75t_R _5687_ (.A(net38),
    .B(_2612_),
    .Y(_2613_));
 OA211x2_ASAP7_75t_R _5688_ (.A1(_2336_),
    .A2(_2353_),
    .B(_2345_),
    .C(_1508_),
    .Y(_2614_));
 INVx2_ASAP7_75t_R _5689_ (.A(_0656_),
    .Y(_2615_));
 OR2x2_ASAP7_75t_R _5690_ (.A(_2615_),
    .B(net229),
    .Y(_2616_));
 OA221x2_ASAP7_75t_R _5691_ (.A1(net38),
    .A2(_2383_),
    .B1(_2613_),
    .B2(_2614_),
    .C(_2616_),
    .Y(_2617_));
 XOR2x2_ASAP7_75t_R _5692_ (.A(_0835_),
    .B(_0660_),
    .Y(_2618_));
 AND4x2_ASAP7_75t_R _5693_ (.A(_2530_),
    .B(_1927_),
    .C(_1855_),
    .D(_2618_),
    .Y(_2619_));
 AO21x2_ASAP7_75t_R _5694_ (.A1(net219),
    .A2(_2617_),
    .B(_2619_),
    .Y(_2620_));
 AND5x2_ASAP7_75t_R _5695_ (.A(net236),
    .B(_2588_),
    .C(_2602_),
    .D(_2611_),
    .E(_2620_),
    .Y(_2621_));
 XNOR2x2_ASAP7_75t_R _5696_ (.A(_0335_),
    .B(_0839_),
    .Y(_2622_));
 INVx2_ASAP7_75t_R _5697_ (.A(_0340_),
    .Y(_2623_));
 XOR2x2_ASAP7_75t_R _5698_ (.A(_0339_),
    .B(_0841_),
    .Y(_2624_));
 NOR2x2_ASAP7_75t_R _5699_ (.A(_2623_),
    .B(_2624_),
    .Y(_2625_));
 AND3x2_ASAP7_75t_R _5700_ (.A(_0336_),
    .B(_2622_),
    .C(_2625_),
    .Y(_2626_));
 XOR2x2_ASAP7_75t_R _5701_ (.A(_0337_),
    .B(_0840_),
    .Y(_2627_));
 INVx2_ASAP7_75t_R _5702_ (.A(_2627_),
    .Y(_2628_));
 AND2x2_ASAP7_75t_R _5703_ (.A(_0338_),
    .B(_2628_),
    .Y(_2629_));
 XOR2x2_ASAP7_75t_R _5704_ (.A(_0333_),
    .B(_0838_),
    .Y(_2630_));
 INVx2_ASAP7_75t_R _5705_ (.A(_2630_),
    .Y(_2631_));
 AND3x2_ASAP7_75t_R _5706_ (.A(_0334_),
    .B(_3709_),
    .C(_2631_),
    .Y(_2632_));
 XOR2x2_ASAP7_75t_R _5707_ (.A(_0665_),
    .B(_0842_),
    .Y(_2633_));
 AND2x2_ASAP7_75t_R _5708_ (.A(_2568_),
    .B(_2633_),
    .Y(_2634_));
 AND3x2_ASAP7_75t_R _5709_ (.A(_2629_),
    .B(_2632_),
    .C(_2634_),
    .Y(_2635_));
 AND3x2_ASAP7_75t_R _5710_ (.A(_1877_),
    .B(_2626_),
    .C(_2635_),
    .Y(_2636_));
 OR2x2_ASAP7_75t_R _5711_ (.A(_2621_),
    .B(_2636_),
    .Y(_3689_));
 XOR2x2_ASAP7_75t_R _5712_ (.A(_0828_),
    .B(_0658_),
    .Y(_2637_));
 OR2x2_ASAP7_75t_R _5713_ (.A(_1598_),
    .B(_2637_),
    .Y(_2638_));
 OR3x2_ASAP7_75t_R _5714_ (.A(_0019_),
    .B(_1849_),
    .C(_1841_),
    .Y(_2639_));
 OR3x2_ASAP7_75t_R _5715_ (.A(_0018_),
    .B(_1842_),
    .C(_1848_),
    .Y(_2640_));
 OR5x2_ASAP7_75t_R _5716_ (.A(_1853_),
    .B(_1621_),
    .C(_1838_),
    .D(_2639_),
    .E(_2640_),
    .Y(_2641_));
 AO211x2_ASAP7_75t_R _5717_ (.A1(_0733_),
    .A2(_2641_),
    .B(_2511_),
    .C(net229),
    .Y(_2642_));
 OA21x2_ASAP7_75t_R _5718_ (.A1(net226),
    .A2(_2638_),
    .B(_2642_),
    .Y(_2643_));
 OA211x2_ASAP7_75t_R _5719_ (.A1(_1677_),
    .A2(_2512_),
    .B(_2528_),
    .C(_2643_),
    .Y(_2644_));
 XOR2x2_ASAP7_75t_R _5720_ (.A(_0663_),
    .B(_2643_),
    .Y(_2645_));
 AND3x2_ASAP7_75t_R _5721_ (.A(_0664_),
    .B(_1877_),
    .C(_2645_),
    .Y(_2646_));
 AO21x2_ASAP7_75t_R _5722_ (.A1(net222),
    .A2(_2644_),
    .B(_2646_),
    .Y(_2647_));
 AND2x2_ASAP7_75t_R _5723_ (.A(_3689_),
    .B(_2647_),
    .Y(_3685_));
 INVx2_ASAP7_75t_R _5724_ (.A(_0843_),
    .Y(_2648_));
 AND2x2_ASAP7_75t_R _5725_ (.A(_2648_),
    .B(_1877_),
    .Y(_2649_));
 INVx2_ASAP7_75t_R _5726_ (.A(_0836_),
    .Y(_2650_));
 AND2x2_ASAP7_75t_R _5727_ (.A(_2650_),
    .B(_1927_),
    .Y(_2651_));
 OR2x2_ASAP7_75t_R _5728_ (.A(_0283_),
    .B(net229),
    .Y(_2652_));
 AO21x2_ASAP7_75t_R _5729_ (.A1(_1855_),
    .A2(_2651_),
    .B(_2652_),
    .Y(_2653_));
 TAPCELL_ASAP7_75t_R PHY_52 ();
 INVx2_ASAP7_75t_R _5731_ (.A(_0283_),
    .Y(_2655_));
 AND2x2_ASAP7_75t_R _5732_ (.A(_2655_),
    .B(net39),
    .Y(_2656_));
 OR4x2_ASAP7_75t_R _5733_ (.A(_0836_),
    .B(_1598_),
    .C(net226),
    .D(_2656_),
    .Y(_2657_));
 TAPCELL_ASAP7_75t_R PHY_51 ();
 AND2x2_ASAP7_75t_R _5735_ (.A(_2653_),
    .B(_2657_),
    .Y(_2659_));
 AND2x2_ASAP7_75t_R _5736_ (.A(_0846_),
    .B(net180),
    .Y(_2660_));
 XNOR2x2_ASAP7_75t_R _5737_ (.A(_2659_),
    .B(_2660_),
    .Y(_2661_));
 XNOR2x2_ASAP7_75t_R _5738_ (.A(_2649_),
    .B(_2661_),
    .Y(_3683_));
 AND3x2_ASAP7_75t_R _5739_ (.A(_0844_),
    .B(_1956_),
    .C(_1961_),
    .Y(_2662_));
 AO21x2_ASAP7_75t_R _5740_ (.A1(net222),
    .A2(_2543_),
    .B(_2662_),
    .Y(_3684_));
 AND2x2_ASAP7_75t_R _5741_ (.A(_0345_),
    .B(net180),
    .Y(_2663_));
 AO21x2_ASAP7_75t_R _5742_ (.A1(net162),
    .A2(_3684_),
    .B(_2663_),
    .Y(_3686_));
 AND2x2_ASAP7_75t_R _5743_ (.A(net228),
    .B(_2529_),
    .Y(_2664_));
 AO21x2_ASAP7_75t_R _5744_ (.A1(_0664_),
    .A2(_1877_),
    .B(_2664_),
    .Y(_3688_));
 AND2x2_ASAP7_75t_R _5745_ (.A(_0348_),
    .B(net180),
    .Y(_2665_));
 AO21x2_ASAP7_75t_R _5746_ (.A1(net162),
    .A2(_3688_),
    .B(_2665_),
    .Y(_3690_));
 OR2x2_ASAP7_75t_R _5747_ (.A(_1877_),
    .B(_2620_),
    .Y(_2666_));
 OA211x2_ASAP7_75t_R _5748_ (.A1(net228),
    .A2(_2634_),
    .B(_2666_),
    .C(_3709_),
    .Y(_2667_));
 TAPCELL_ASAP7_75t_R PHY_50 ();
 AND2x2_ASAP7_75t_R _5750_ (.A(net222),
    .B(_2588_),
    .Y(_2668_));
 AO32x2_ASAP7_75t_R _5751_ (.A1(_1877_),
    .A2(_2629_),
    .A3(_2626_),
    .B1(_2602_),
    .B2(_2668_),
    .Y(_2669_));
 AND2x2_ASAP7_75t_R _5752_ (.A(_2667_),
    .B(_2669_),
    .Y(_3693_));
 AND2x2_ASAP7_75t_R _5753_ (.A(_0852_),
    .B(net180),
    .Y(_2670_));
 AND2x2_ASAP7_75t_R _5754_ (.A(net223),
    .B(_2603_),
    .Y(_2671_));
 AO21x2_ASAP7_75t_R _5755_ (.A1(net229),
    .A2(_3337_),
    .B(_2671_),
    .Y(_3662_));
 OR2x2_ASAP7_75t_R _5756_ (.A(_1677_),
    .B(_3662_),
    .Y(_2672_));
 OA21x2_ASAP7_75t_R _5757_ (.A1(net219),
    .A2(_2608_),
    .B(_2672_),
    .Y(_3672_));
 AND2x2_ASAP7_75t_R _5758_ (.A(_1877_),
    .B(_2630_),
    .Y(_2673_));
 AO21x2_ASAP7_75t_R _5759_ (.A1(net222),
    .A2(_3672_),
    .B(_2673_),
    .Y(_2674_));
 XNOR2x2_ASAP7_75t_R _5760_ (.A(_2670_),
    .B(_2674_),
    .Y(_3691_));
 AND2x2_ASAP7_75t_R _5761_ (.A(net162),
    .B(_3692_),
    .Y(_2675_));
 AND2x2_ASAP7_75t_R _5762_ (.A(_0353_),
    .B(net180),
    .Y(_2676_));
 OR2x2_ASAP7_75t_R _5763_ (.A(_2675_),
    .B(_2676_),
    .Y(_3694_));
 AND2x2_ASAP7_75t_R _5764_ (.A(_0854_),
    .B(net180),
    .Y(_2677_));
 INVx2_ASAP7_75t_R _5765_ (.A(_2591_),
    .Y(_2678_));
 OR2x2_ASAP7_75t_R _5766_ (.A(_1677_),
    .B(_2595_),
    .Y(_2679_));
 OA21x2_ASAP7_75t_R _5767_ (.A1(net219),
    .A2(_2678_),
    .B(_2679_),
    .Y(_3673_));
 NOR2x2_ASAP7_75t_R _5768_ (.A(net222),
    .B(_2622_),
    .Y(_2680_));
 AO21x2_ASAP7_75t_R _5769_ (.A1(net222),
    .A2(_3673_),
    .B(_2680_),
    .Y(_2681_));
 XNOR2x2_ASAP7_75t_R _5770_ (.A(_2677_),
    .B(_2681_),
    .Y(_3695_));
 AND2x2_ASAP7_75t_R _5771_ (.A(net162),
    .B(_3696_),
    .Y(_2682_));
 AND2x2_ASAP7_75t_R _5772_ (.A(_0358_),
    .B(net180),
    .Y(_2683_));
 OR2x2_ASAP7_75t_R _5773_ (.A(_2682_),
    .B(_2683_),
    .Y(_3698_));
 AO221x2_ASAP7_75t_R _5774_ (.A1(_1956_),
    .A2(_1961_),
    .B1(_2590_),
    .B2(_1677_),
    .C(_2601_),
    .Y(_2684_));
 OA211x2_ASAP7_75t_R _5775_ (.A1(net222),
    .A2(_2625_),
    .B(_2667_),
    .C(_2684_),
    .Y(_3701_));
 AND2x2_ASAP7_75t_R _5776_ (.A(_0856_),
    .B(net180),
    .Y(_2685_));
 OR2x2_ASAP7_75t_R _5777_ (.A(_1677_),
    .B(_2583_),
    .Y(_2686_));
 OA21x2_ASAP7_75t_R _5778_ (.A1(net219),
    .A2(_2585_),
    .B(_2686_),
    .Y(_3674_));
 AND2x2_ASAP7_75t_R _5779_ (.A(_1877_),
    .B(_2627_),
    .Y(_2687_));
 AO21x2_ASAP7_75t_R _5780_ (.A1(net222),
    .A2(_3674_),
    .B(_2687_),
    .Y(_2688_));
 XNOR2x2_ASAP7_75t_R _5781_ (.A(_2685_),
    .B(_2688_),
    .Y(_3699_));
 AND2x2_ASAP7_75t_R _5782_ (.A(net162),
    .B(_3700_),
    .Y(_2689_));
 AND2x2_ASAP7_75t_R _5783_ (.A(_0362_),
    .B(net180),
    .Y(_2690_));
 OR2x2_ASAP7_75t_R _5784_ (.A(_2689_),
    .B(_2690_),
    .Y(_3702_));
 AND2x2_ASAP7_75t_R _5785_ (.A(_0858_),
    .B(net180),
    .Y(_2691_));
 AND2x2_ASAP7_75t_R _5786_ (.A(net233),
    .B(_2597_),
    .Y(_2692_));
 AO21x2_ASAP7_75t_R _5787_ (.A1(net229),
    .A2(_2315_),
    .B(_2692_),
    .Y(_3665_));
 AND2x2_ASAP7_75t_R _5788_ (.A(net219),
    .B(_3665_),
    .Y(_2693_));
 AO21x2_ASAP7_75t_R _5789_ (.A1(_1677_),
    .A2(_2589_),
    .B(_2693_),
    .Y(_3675_));
 OR2x2_ASAP7_75t_R _5790_ (.A(net222),
    .B(_2624_),
    .Y(_2694_));
 OA21x2_ASAP7_75t_R _5791_ (.A1(_1877_),
    .A2(_3675_),
    .B(_2694_),
    .Y(_2695_));
 XNOR2x2_ASAP7_75t_R _5792_ (.A(_2691_),
    .B(_2695_),
    .Y(_3703_));
 AND2x2_ASAP7_75t_R _5793_ (.A(net162),
    .B(_3704_),
    .Y(_2696_));
 AND2x2_ASAP7_75t_R _5794_ (.A(_0367_),
    .B(net180),
    .Y(_2697_));
 OR2x2_ASAP7_75t_R _5795_ (.A(_2696_),
    .B(_2697_),
    .Y(_3706_));
 AND2x2_ASAP7_75t_R _5796_ (.A(_0860_),
    .B(net180),
    .Y(_2698_));
 XNOR2x2_ASAP7_75t_R _5797_ (.A(_0835_),
    .B(_0660_),
    .Y(_2699_));
 NOR2x2_ASAP7_75t_R _5798_ (.A(_2613_),
    .B(_2614_),
    .Y(_3666_));
 OR2x2_ASAP7_75t_R _5799_ (.A(_1677_),
    .B(_3666_),
    .Y(_2700_));
 OA21x2_ASAP7_75t_R _5800_ (.A1(net221),
    .A2(_2699_),
    .B(_2700_),
    .Y(_3676_));
 AND2x2_ASAP7_75t_R _5801_ (.A(net228),
    .B(_3676_),
    .Y(_2701_));
 INVx2_ASAP7_75t_R _5802_ (.A(_2701_),
    .Y(_2702_));
 OA21x2_ASAP7_75t_R _5803_ (.A1(net228),
    .A2(_2633_),
    .B(_2702_),
    .Y(_2703_));
 XOR2x2_ASAP7_75t_R _5804_ (.A(_2698_),
    .B(_2703_),
    .Y(_3707_));
 AND2x2_ASAP7_75t_R _5805_ (.A(net162),
    .B(_3708_),
    .Y(_2704_));
 AND2x2_ASAP7_75t_R _5806_ (.A(_0371_),
    .B(net180),
    .Y(_2705_));
 OR2x2_ASAP7_75t_R _5807_ (.A(_2704_),
    .B(_2705_),
    .Y(_3710_));
 INVx2_ASAP7_75t_R _5808_ (.A(_3721_),
    .Y(_3376_));
 OA21x2_ASAP7_75t_R _5809_ (.A1(_0374_),
    .A2(_3376_),
    .B(_0372_),
    .Y(_2706_));
 OA21x2_ASAP7_75t_R _5810_ (.A1(_0859_),
    .A2(_2706_),
    .B(_0370_),
    .Y(_3381_));
 OA21x2_ASAP7_75t_R _5811_ (.A1(_0369_),
    .A2(_3381_),
    .B(_0368_),
    .Y(_2707_));
 OA21x2_ASAP7_75t_R _5812_ (.A1(_0857_),
    .A2(_2707_),
    .B(_0365_),
    .Y(_3384_));
 OA21x2_ASAP7_75t_R _5813_ (.A1(_0364_),
    .A2(_3384_),
    .B(_0363_),
    .Y(_2708_));
 OA21x2_ASAP7_75t_R _5814_ (.A1(_0855_),
    .A2(_2708_),
    .B(_0361_),
    .Y(_3387_));
 OA211x2_ASAP7_75t_R _5815_ (.A1(_0855_),
    .A2(_2708_),
    .B(_0359_),
    .C(_0361_),
    .Y(_2709_));
 AO21x2_ASAP7_75t_R _5816_ (.A1(_0359_),
    .A2(_0360_),
    .B(_0853_),
    .Y(_2710_));
 AND3x2_ASAP7_75t_R _5817_ (.A(_0354_),
    .B(_0357_),
    .C(_0850_),
    .Y(_2711_));
 OA21x2_ASAP7_75t_R _5818_ (.A1(_2709_),
    .A2(_2710_),
    .B(_2711_),
    .Y(_2712_));
 AND2x2_ASAP7_75t_R _5819_ (.A(_0354_),
    .B(_0355_),
    .Y(_2713_));
 OA21x2_ASAP7_75t_R _5820_ (.A1(_0851_),
    .A2(_2713_),
    .B(_0850_),
    .Y(_2714_));
 OR2x2_ASAP7_75t_R _5821_ (.A(_2712_),
    .B(_2714_),
    .Y(_3393_));
 OA21x2_ASAP7_75t_R _5822_ (.A1(_0351_),
    .A2(_3393_),
    .B(_0349_),
    .Y(_2715_));
 OA21x2_ASAP7_75t_R _5823_ (.A1(_0848_),
    .A2(_2715_),
    .B(_0847_),
    .Y(_3396_));
 OR2x2_ASAP7_75t_R _5824_ (.A(_0289_),
    .B(_0828_),
    .Y(_2716_));
 OA21x2_ASAP7_75t_R _5825_ (.A1(_0288_),
    .A2(_0828_),
    .B(_0286_),
    .Y(_2717_));
 OA21x2_ASAP7_75t_R _5826_ (.A1(_3314_),
    .A2(_2716_),
    .B(_2717_),
    .Y(_2718_));
 OR4x2_ASAP7_75t_R _5827_ (.A(_0283_),
    .B(net219),
    .C(_2510_),
    .D(_2718_),
    .Y(_2719_));
 INVx2_ASAP7_75t_R _5828_ (.A(_2719_),
    .Y(_3713_));
 OR2x2_ASAP7_75t_R _5829_ (.A(_1877_),
    .B(_2719_),
    .Y(_2720_));
 OA21x2_ASAP7_75t_R _5830_ (.A1(_0379_),
    .A2(net222),
    .B(_2720_),
    .Y(_3716_));
 AND3x2_ASAP7_75t_R _5831_ (.A(net222),
    .B(_2644_),
    .C(_2719_),
    .Y(_2721_));
 AND2x2_ASAP7_75t_R _5832_ (.A(_0378_),
    .B(_0379_),
    .Y(_2722_));
 AND4x2_ASAP7_75t_R _5833_ (.A(_0664_),
    .B(_1877_),
    .C(_2645_),
    .D(_2722_),
    .Y(_2723_));
 NAND3x2_ASAP7_75t_R _5834_ (.B(_2653_),
    .C(_2657_),
    .Y(_2724_),
    .A(_2648_));
 AO21x2_ASAP7_75t_R _5835_ (.A1(_2653_),
    .A2(_2657_),
    .B(_2648_),
    .Y(_2725_));
 AO33x2_ASAP7_75t_R _5836_ (.A1(net222),
    .A2(_2543_),
    .A3(_2659_),
    .B1(_2662_),
    .B2(_2724_),
    .B3(_2725_),
    .Y(_2726_));
 OA221x2_ASAP7_75t_R _5837_ (.A1(_2621_),
    .A2(_2636_),
    .B1(_2721_),
    .B2(_2723_),
    .C(_2726_),
    .Y(_2727_));
 NOR2x2_ASAP7_75t_R _5838_ (.A(net162),
    .B(_2727_),
    .Y(_3357_));
 OR2x2_ASAP7_75t_R _5839_ (.A(_0378_),
    .B(net222),
    .Y(_2728_));
 AND2x2_ASAP7_75t_R _5840_ (.A(_0867_),
    .B(net180),
    .Y(_2729_));
 XOR2x2_ASAP7_75t_R _5841_ (.A(_2728_),
    .B(_2729_),
    .Y(_3715_));
 AND2x2_ASAP7_75t_R _5842_ (.A(_0404_),
    .B(net180),
    .Y(_2730_));
 AO21x2_ASAP7_75t_R _5843_ (.A1(net162),
    .A2(_3716_),
    .B(_2730_),
    .Y(_3371_));
 AO21x2_ASAP7_75t_R _5844_ (.A1(_0847_),
    .A2(_0848_),
    .B(_0347_),
    .Y(_2731_));
 AO21x2_ASAP7_75t_R _5845_ (.A1(_0346_),
    .A2(_2731_),
    .B(_0344_),
    .Y(_2732_));
 AND2x2_ASAP7_75t_R _5846_ (.A(_0407_),
    .B(_2732_),
    .Y(_2733_));
 OR5x2_ASAP7_75t_R _5847_ (.A(_0406_),
    .B(_0351_),
    .C(_2712_),
    .D(_2714_),
    .E(_2733_),
    .Y(_2734_));
 AND3x2_ASAP7_75t_R _5848_ (.A(_0346_),
    .B(_0407_),
    .C(_0847_),
    .Y(_2735_));
 AO221x2_ASAP7_75t_R _5849_ (.A1(_0349_),
    .A2(_2735_),
    .B1(_2732_),
    .B2(_0407_),
    .C(_0406_),
    .Y(_2736_));
 AND3x2_ASAP7_75t_R _5850_ (.A(_0400_),
    .B(_0405_),
    .C(_0402_),
    .Y(_2737_));
 AND3x2_ASAP7_75t_R _5851_ (.A(_0400_),
    .B(_0403_),
    .C(_0402_),
    .Y(_2738_));
 AO21x2_ASAP7_75t_R _5852_ (.A1(_0400_),
    .A2(_0401_),
    .B(_2738_),
    .Y(_2739_));
 AO31x2_ASAP7_75t_R _5853_ (.A1(_2734_),
    .A2(_2736_),
    .A3(_2737_),
    .B(_2739_),
    .Y(_2740_));
 OR3x2_ASAP7_75t_R _5854_ (.A(_0398_),
    .B(_0865_),
    .C(_0866_),
    .Y(_2741_));
 OR2x2_ASAP7_75t_R _5855_ (.A(_0398_),
    .B(_0399_),
    .Y(_2742_));
 AO21x2_ASAP7_75t_R _5856_ (.A1(_0396_),
    .A2(_2742_),
    .B(_0865_),
    .Y(_2743_));
 AND3x2_ASAP7_75t_R _5857_ (.A(_0393_),
    .B(_0391_),
    .C(_0395_),
    .Y(_2744_));
 OA211x2_ASAP7_75t_R _5858_ (.A1(_2740_),
    .A2(_2741_),
    .B(_2743_),
    .C(_2744_),
    .Y(_2745_));
 AND3x2_ASAP7_75t_R _5859_ (.A(_0393_),
    .B(_0391_),
    .C(_0394_),
    .Y(_2746_));
 AO21x2_ASAP7_75t_R _5860_ (.A1(_0391_),
    .A2(_0864_),
    .B(_2746_),
    .Y(_2747_));
 OR2x2_ASAP7_75t_R _5861_ (.A(_2745_),
    .B(_2747_),
    .Y(_3364_));
 OR2x2_ASAP7_75t_R _5862_ (.A(_0387_),
    .B(_0390_),
    .Y(_2748_));
 OA21x2_ASAP7_75t_R _5863_ (.A1(_0388_),
    .A2(_0387_),
    .B(_0863_),
    .Y(_2749_));
 OA31x2_ASAP7_75t_R _5864_ (.A1(_2745_),
    .A2(_2747_),
    .A3(_2748_),
    .B1(_2749_),
    .Y(_3362_));
 OR2x2_ASAP7_75t_R _5865_ (.A(_0384_),
    .B(_0386_),
    .Y(_2750_));
 OA21x2_ASAP7_75t_R _5866_ (.A1(_0385_),
    .A2(_0384_),
    .B(_0862_),
    .Y(_2751_));
 OA21x2_ASAP7_75t_R _5867_ (.A1(_3362_),
    .A2(_2750_),
    .B(_2751_),
    .Y(_3360_));
 OA21x2_ASAP7_75t_R _5868_ (.A1(_0383_),
    .A2(_3360_),
    .B(_0382_),
    .Y(_2752_));
 OA21x2_ASAP7_75t_R _5869_ (.A1(_0381_),
    .A2(_2752_),
    .B(_0861_),
    .Y(_3358_));
 OA21x2_ASAP7_75t_R _5870_ (.A1(_0866_),
    .A2(_2740_),
    .B(_0399_),
    .Y(_3368_));
 AND3x2_ASAP7_75t_R _5871_ (.A(_0405_),
    .B(_2734_),
    .C(_2736_),
    .Y(_2753_));
 OA21x2_ASAP7_75t_R _5872_ (.A1(_0403_),
    .A2(_2753_),
    .B(_0402_),
    .Y(_3370_));
 OA21x2_ASAP7_75t_R _5873_ (.A1(_2709_),
    .A2(_2710_),
    .B(_0357_),
    .Y(_3390_));
 INVx2_ASAP7_75t_R _5874_ (.A(_0515_),
    .Y(net37));
 OR2x4_ASAP7_75t_R _5875_ (.A(net18),
    .B(_0515_),
    .Y(_2754_));
 OR2x2_ASAP7_75t_R _5876_ (.A(_0427_),
    .B(_2754_),
    .Y(_2755_));
 NAND2x2_ASAP7_75t_R _5877_ (.A(net17),
    .B(_2755_),
    .Y(_2756_));
 INVx6_ASAP7_75t_R _5878_ (.A(_2756_),
    .Y(net20));
 TAPCELL_ASAP7_75t_R PHY_49 ();
 BUFx4_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 INVx2_ASAP7_75t_R _5881_ (.A(_0516_),
    .Y(\__in_sample_reg[14] ));
 INVx2_ASAP7_75t_R _5882_ (.A(_0517_),
    .Y(\__in_sample_reg[13] ));
 INVx2_ASAP7_75t_R _5883_ (.A(_0518_),
    .Y(\__in_sample_reg[12] ));
 INVx2_ASAP7_75t_R _5884_ (.A(_0519_),
    .Y(\__in_sample_reg[11] ));
 INVx2_ASAP7_75t_R _5885_ (.A(_0520_),
    .Y(\__in_sample_reg[10] ));
 INVx2_ASAP7_75t_R _5886_ (.A(_0521_),
    .Y(\__in_sample_reg[9] ));
 INVx2_ASAP7_75t_R _5887_ (.A(_0522_),
    .Y(\__in_sample_reg[8] ));
 INVx2_ASAP7_75t_R _5888_ (.A(_0523_),
    .Y(\__in_sample_reg[7] ));
 INVx2_ASAP7_75t_R _5889_ (.A(_0524_),
    .Y(\__in_sample_reg[6] ));
 INVx2_ASAP7_75t_R _5890_ (.A(_0525_),
    .Y(\__in_sample_reg[5] ));
 INVx2_ASAP7_75t_R _5891_ (.A(_3129_),
    .Y(\__in_sample_reg[4] ));
 INVx2_ASAP7_75t_R _5892_ (.A(_0526_),
    .Y(\__in_sample_reg[3] ));
 INVx2_ASAP7_75t_R _5893_ (.A(_0527_),
    .Y(\__in_sample_reg[2] ));
 INVx2_ASAP7_75t_R _5894_ (.A(_0528_),
    .Y(\__in_sample_reg[1] ));
 INVx2_ASAP7_75t_R _5895_ (.A(_0530_),
    .Y(\__st_3[29] ));
 INVx2_ASAP7_75t_R _5896_ (.A(_3359_),
    .Y(\__st_3[28] ));
 INVx2_ASAP7_75t_R _5897_ (.A(_0531_),
    .Y(\__st_3[27] ));
 INVx2_ASAP7_75t_R _5898_ (.A(_3361_),
    .Y(\__st_3[26] ));
 INVx2_ASAP7_75t_R _5899_ (.A(_0532_),
    .Y(\__st_3[25] ));
 INVx2_ASAP7_75t_R _5900_ (.A(_3363_),
    .Y(\__st_3[24] ));
 INVx2_ASAP7_75t_R _5901_ (.A(_0533_),
    .Y(\__st_3[23] ));
 INVx2_ASAP7_75t_R _5902_ (.A(_0534_),
    .Y(\__st_3[22] ));
 INVx2_ASAP7_75t_R _5903_ (.A(_0535_),
    .Y(\__st_3[21] ));
 INVx2_ASAP7_75t_R _5904_ (.A(_3367_),
    .Y(\__st_3[20] ));
 INVx2_ASAP7_75t_R _5905_ (.A(_0536_),
    .Y(\__st_3[19] ));
 INVx2_ASAP7_75t_R _5906_ (.A(_3369_),
    .Y(\__st_3[18] ));
 INVx2_ASAP7_75t_R _5907_ (.A(_0537_),
    .Y(\__st_3[17] ));
 INVx2_ASAP7_75t_R _5908_ (.A(_0538_),
    .Y(\__st_3[16] ));
 INVx2_ASAP7_75t_R _5909_ (.A(_0539_),
    .Y(net27));
 INVx2_ASAP7_75t_R _5910_ (.A(_3394_),
    .Y(net26));
 INVx2_ASAP7_75t_R _5911_ (.A(_0540_),
    .Y(net25));
 INVx2_ASAP7_75t_R _5912_ (.A(_3391_),
    .Y(net24));
 INVx2_ASAP7_75t_R _5913_ (.A(_0541_),
    .Y(net23));
 INVx2_ASAP7_75t_R _5914_ (.A(_3388_),
    .Y(net22));
 INVx2_ASAP7_75t_R _5915_ (.A(_0542_),
    .Y(net36));
 INVx2_ASAP7_75t_R _5916_ (.A(_3385_),
    .Y(net35));
 INVx2_ASAP7_75t_R _5917_ (.A(_0543_),
    .Y(net34));
 INVx2_ASAP7_75t_R _5918_ (.A(_3382_),
    .Y(net33));
 INVx2_ASAP7_75t_R _5919_ (.A(_0544_),
    .Y(net32));
 INVx2_ASAP7_75t_R _5920_ (.A(_3379_),
    .Y(net31));
 INVx2_ASAP7_75t_R _5921_ (.A(_0545_),
    .Y(net30));
 INVx2_ASAP7_75t_R _5922_ (.A(_3377_),
    .Y(net29));
 INVx2_ASAP7_75t_R _5923_ (.A(_3373_),
    .Y(net28));
 INVx2_ASAP7_75t_R _5924_ (.A(_3718_),
    .Y(net21));
 INVx2_ASAP7_75t_R _5925_ (.A(_3411_),
    .Y(\__st_1[29] ));
 INVx2_ASAP7_75t_R _5926_ (.A(_3141_),
    .Y(\__st_1[28] ));
 INVx2_ASAP7_75t_R _5927_ (.A(_3412_),
    .Y(\__st_1[27] ));
 INVx2_ASAP7_75t_R _5928_ (.A(_3143_),
    .Y(\__st_1[26] ));
 INVx2_ASAP7_75t_R _5929_ (.A(_3413_),
    .Y(\__st_1[25] ));
 INVx2_ASAP7_75t_R _5930_ (.A(_3258_),
    .Y(\__st_1[24] ));
 INVx2_ASAP7_75t_R _5931_ (.A(_3414_),
    .Y(\__st_1[23] ));
 INVx3_ASAP7_75t_R _5932_ (.A(_3415_),
    .Y(\__st_1[22] ));
 INVx2_ASAP7_75t_R _5933_ (.A(_3416_),
    .Y(\__st_1[21] ));
 INVx2_ASAP7_75t_R _5934_ (.A(_3262_),
    .Y(\__st_1[20] ));
 INVx2_ASAP7_75t_R _5935_ (.A(_3417_),
    .Y(\__st_1[19] ));
 INVx3_ASAP7_75t_R _5936_ (.A(_3418_),
    .Y(\__st_1[18] ));
 INVx2_ASAP7_75t_R _5937_ (.A(_3419_),
    .Y(\__st_1[17] ));
 INVx2_ASAP7_75t_R _5938_ (.A(_3265_),
    .Y(\__st_1[16] ));
 INVx2_ASAP7_75t_R _5939_ (.A(_3420_),
    .Y(\__st_1[15] ));
 INVx2_ASAP7_75t_R _5940_ (.A(_3131_),
    .Y(\__st_1[14] ));
 INVx2_ASAP7_75t_R _5941_ (.A(_3421_),
    .Y(\__st_1[13] ));
 INVx2_ASAP7_75t_R _5942_ (.A(_3133_),
    .Y(\__st_1[12] ));
 INVx2_ASAP7_75t_R _5943_ (.A(_3422_),
    .Y(\__st_1[11] ));
 INVx2_ASAP7_75t_R _5944_ (.A(_3135_),
    .Y(\__st_1[10] ));
 INVx2_ASAP7_75t_R _5945_ (.A(_3423_),
    .Y(\__st_1[9] ));
 INVx2_ASAP7_75t_R _5946_ (.A(_3137_),
    .Y(\__st_1[8] ));
 INVx2_ASAP7_75t_R _5947_ (.A(_3424_),
    .Y(\__st_1[7] ));
 INVx2_ASAP7_75t_R _5948_ (.A(_3127_),
    .Y(\__st_1[6] ));
 INVx2_ASAP7_75t_R _5949_ (.A(_3425_),
    .Y(\__st_1[5] ));
 INVx2_ASAP7_75t_R _5950_ (.A(_3272_),
    .Y(\__st_1[4] ));
 INVx2_ASAP7_75t_R _5951_ (.A(_3426_),
    .Y(\__st_1[3] ));
 INVx2_ASAP7_75t_R _5952_ (.A(_3126_),
    .Y(\__st_1[2] ));
 INVx2_ASAP7_75t_R _5953_ (.A(_3584_),
    .Y(\__st_1[0] ));
 INVx2_ASAP7_75t_R _5954_ (.A(_2459_),
    .Y(_3308_));
 INVx2_ASAP7_75t_R _5955_ (.A(_3616_),
    .Y(_3266_));
 INVx2_ASAP7_75t_R _5956_ (.A(_0240_),
    .Y(_2758_));
 OR2x2_ASAP7_75t_R _5957_ (.A(_2758_),
    .B(net162),
    .Y(_2759_));
 OA21x2_ASAP7_75t_R _5958_ (.A1(net180),
    .A2(_2002_),
    .B(_2759_),
    .Y(_3268_));
 NOR2x2_ASAP7_75t_R _5959_ (.A(_2131_),
    .B(_2132_),
    .Y(_3271_));
 NOR2x2_ASAP7_75t_R _5960_ (.A(_2122_),
    .B(_2123_),
    .Y(_3273_));
 NOR2x2_ASAP7_75t_R _5961_ (.A(_2118_),
    .B(_2119_),
    .Y(_3275_));
 NOR2x2_ASAP7_75t_R _5962_ (.A(_2101_),
    .B(_2102_),
    .Y(_3277_));
 INVx2_ASAP7_75t_R _5963_ (.A(_3627_),
    .Y(_3279_));
 INVx2_ASAP7_75t_R _5964_ (.A(_3623_),
    .Y(_3281_));
 INVx2_ASAP7_75t_R _5965_ (.A(_0375_),
    .Y(_2760_));
 OR2x2_ASAP7_75t_R _5966_ (.A(_2760_),
    .B(net162),
    .Y(_2761_));
 OA21x2_ASAP7_75t_R _5967_ (.A1(net180),
    .A2(_2573_),
    .B(_2761_),
    .Y(_3374_));
 NOR2x2_ASAP7_75t_R _5968_ (.A(_2704_),
    .B(_2705_),
    .Y(_3378_));
 NOR2x2_ASAP7_75t_R _5969_ (.A(_2696_),
    .B(_2697_),
    .Y(_3380_));
 NOR2x2_ASAP7_75t_R _5970_ (.A(_2689_),
    .B(_2690_),
    .Y(_3383_));
 NOR2x2_ASAP7_75t_R _5971_ (.A(_2682_),
    .B(_2683_),
    .Y(_3386_));
 NOR2x2_ASAP7_75t_R _5972_ (.A(_2675_),
    .B(_2676_),
    .Y(_3389_));
 INVx2_ASAP7_75t_R _5973_ (.A(_3690_),
    .Y(_3392_));
 INVx2_ASAP7_75t_R _5974_ (.A(_3686_),
    .Y(_3395_));
 OR2x2_ASAP7_75t_R _5975_ (.A(_3206_),
    .B(_0995_),
    .Y(_3400_));
 OR2x2_ASAP7_75t_R _5976_ (.A(_1151_),
    .B(_1153_),
    .Y(_2762_));
 INVx2_ASAP7_75t_R _5977_ (.A(_2762_),
    .Y(_3134_));
 INVx2_ASAP7_75t_R _5978_ (.A(_1148_),
    .Y(_3138_));
 OR2x2_ASAP7_75t_R _5979_ (.A(_0392_),
    .B(_0408_),
    .Y(_2763_));
 OR2x2_ASAP7_75t_R _5980_ (.A(_0410_),
    .B(_2763_),
    .Y(_2764_));
 OA222x2_ASAP7_75t_R _5981_ (.A1(_0397_),
    .A2(_0392_),
    .B1(_0409_),
    .B2(_2763_),
    .C1(_2764_),
    .C2(_1170_),
    .Y(_2765_));
 AND3x2_ASAP7_75t_R _5982_ (.A(_0377_),
    .B(_0373_),
    .C(_0389_),
    .Y(_2766_));
 AND3x2_ASAP7_75t_R _5983_ (.A(_0377_),
    .B(_0373_),
    .C(_0380_),
    .Y(_2767_));
 AO221x2_ASAP7_75t_R _5984_ (.A1(_0376_),
    .A2(_0373_),
    .B1(_2765_),
    .B2(_2766_),
    .C(_2767_),
    .Y(_2768_));
 INVx2_ASAP7_75t_R _5985_ (.A(_2768_),
    .Y(_3142_));
 AND2x2_ASAP7_75t_R _5986_ (.A(_0717_),
    .B(net162),
    .Y(_2769_));
 AO21x2_ASAP7_75t_R _5987_ (.A1(_3479_),
    .A2(net209),
    .B(_2769_),
    .Y(_3495_));
 AND2x2_ASAP7_75t_R _5988_ (.A(_0722_),
    .B(net195),
    .Y(_2770_));
 AO21x2_ASAP7_75t_R _5989_ (.A1(_3485_),
    .A2(net209),
    .B(_2770_),
    .Y(_3501_));
 OR2x2_ASAP7_75t_R _5990_ (.A(_1538_),
    .B(_1539_),
    .Y(_3507_));
 AND2x2_ASAP7_75t_R _5991_ (.A(_0728_),
    .B(net195),
    .Y(_2771_));
 AO21x2_ASAP7_75t_R _5992_ (.A1(_3493_),
    .A2(net209),
    .B(_2771_),
    .Y(_3509_));
 OR2x2_ASAP7_75t_R _5993_ (.A(_3155_),
    .B(net39),
    .Y(_2772_));
 OA21x2_ASAP7_75t_R _5994_ (.A1(_1607_),
    .A2(_1508_),
    .B(_2772_),
    .Y(_3553_));
 INVx2_ASAP7_75t_R _5995_ (.A(_1703_),
    .Y(_3190_));
 INVx2_ASAP7_75t_R _5996_ (.A(_0013_),
    .Y(_2773_));
 OR2x2_ASAP7_75t_R _5997_ (.A(net233),
    .B(_3495_),
    .Y(_2774_));
 OA21x2_ASAP7_75t_R _5998_ (.A1(_2773_),
    .A2(_1508_),
    .B(_2774_),
    .Y(_3560_));
 INVx2_ASAP7_75t_R _5999_ (.A(_0014_),
    .Y(_2775_));
 OR2x2_ASAP7_75t_R _6000_ (.A(_3497_),
    .B(net39),
    .Y(_2776_));
 OA21x2_ASAP7_75t_R _6001_ (.A1(_2775_),
    .A2(_1508_),
    .B(_2776_),
    .Y(_3562_));
 OR2x2_ASAP7_75t_R _6002_ (.A(_3499_),
    .B(_1507_),
    .Y(_2777_));
 OA21x2_ASAP7_75t_R _6003_ (.A1(_1666_),
    .A2(_1508_),
    .B(_2777_),
    .Y(_3564_));
 OR2x2_ASAP7_75t_R _6004_ (.A(_1507_),
    .B(_3501_),
    .Y(_2778_));
 OA21x2_ASAP7_75t_R _6005_ (.A1(_1667_),
    .A2(_1508_),
    .B(_2778_),
    .Y(_3566_));
 INVx2_ASAP7_75t_R _6006_ (.A(_0017_),
    .Y(_2779_));
 OR2x2_ASAP7_75t_R _6007_ (.A(_1507_),
    .B(_1532_),
    .Y(_2780_));
 OA21x2_ASAP7_75t_R _6008_ (.A1(_2779_),
    .A2(_1508_),
    .B(_2780_),
    .Y(_3568_));
 OR2x2_ASAP7_75t_R _6009_ (.A(net39),
    .B(_3505_),
    .Y(_2781_));
 OA21x2_ASAP7_75t_R _6010_ (.A1(_1653_),
    .A2(_1508_),
    .B(_2781_),
    .Y(_3570_));
 OR2x2_ASAP7_75t_R _6011_ (.A(_3507_),
    .B(net39),
    .Y(_2782_));
 OA21x2_ASAP7_75t_R _6012_ (.A1(_1652_),
    .A2(_1508_),
    .B(_2782_),
    .Y(_3572_));
 INVx2_ASAP7_75t_R _6013_ (.A(_0020_),
    .Y(_2783_));
 OR2x2_ASAP7_75t_R _6014_ (.A(net39),
    .B(_3509_),
    .Y(_2784_));
 OA21x2_ASAP7_75t_R _6015_ (.A1(_2783_),
    .A2(_1508_),
    .B(_2784_),
    .Y(_3574_));
 NAND2x2_ASAP7_75t_R _6016_ (.A(_0513_),
    .B(_1872_),
    .Y(_3205_));
 CKINVDCx5p33_ASAP7_75t_R _6017_ (.A(_1363_),
    .Y(_3191_));
 AO32x2_ASAP7_75t_R _6018_ (.A1(net236),
    .A2(_1972_),
    .A3(_1975_),
    .B1(_2093_),
    .B2(_2048_),
    .Y(_2785_));
 AND2x2_ASAP7_75t_R _6019_ (.A(_3626_),
    .B(_2785_),
    .Y(_3622_));
 OR2x2_ASAP7_75t_R _6020_ (.A(_1906_),
    .B(_2125_),
    .Y(_2786_));
 OR3x2_ASAP7_75t_R _6021_ (.A(_0604_),
    .B(net219),
    .C(_2026_),
    .Y(_2787_));
 OA21x2_ASAP7_75t_R _6022_ (.A1(_1677_),
    .A2(_2786_),
    .B(_2787_),
    .Y(_2788_));
 NAND2x2_ASAP7_75t_R _6023_ (.A(_1864_),
    .B(_2788_),
    .Y(_2789_));
 OA211x2_ASAP7_75t_R _6024_ (.A1(net236),
    .A2(_2107_),
    .B(_2789_),
    .C(_3642_),
    .Y(_3638_));
 NAND2x2_ASAP7_75t_R _6025_ (.A(_0254_),
    .B(_2173_),
    .Y(_3291_));
 NAND2x2_ASAP7_75t_R _6026_ (.A(_0259_),
    .B(_2187_),
    .Y(_3650_));
 OR2x2_ASAP7_75t_R _6027_ (.A(_0565_),
    .B(_2185_),
    .Y(_3656_));
 OR2x2_ASAP7_75t_R _6028_ (.A(_2575_),
    .B(_2580_),
    .Y(_3719_));
 OR2x2_ASAP7_75t_R _6029_ (.A(_0555_),
    .B(_0995_),
    .Y(_3398_));
 INVx2_ASAP7_75t_R _6030_ (.A(_1183_),
    .Y(_3175_));
 INVx2_ASAP7_75t_R _6031_ (.A(_3430_),
    .Y(_3431_));
 INVx2_ASAP7_75t_R _6032_ (.A(_1238_),
    .Y(_3172_));
 INVx2_ASAP7_75t_R _6033_ (.A(_1146_),
    .Y(_3128_));
 INVx2_ASAP7_75t_R _6034_ (.A(_3437_),
    .Y(_3438_));
 INVx2_ASAP7_75t_R _6035_ (.A(_1293_),
    .Y(_3166_));
 INVx2_ASAP7_75t_R _6036_ (.A(_3446_),
    .Y(_3447_));
 INVx2_ASAP7_75t_R _6037_ (.A(_1338_),
    .Y(_3169_));
 OA21x2_ASAP7_75t_R _6038_ (.A1(_0435_),
    .A2(_2762_),
    .B(_0434_),
    .Y(_2790_));
 OA21x2_ASAP7_75t_R _6039_ (.A1(_0702_),
    .A2(_2790_),
    .B(_0433_),
    .Y(_2791_));
 INVx2_ASAP7_75t_R _6040_ (.A(_2791_),
    .Y(_3132_));
 OA21x2_ASAP7_75t_R _6041_ (.A1(_0704_),
    .A2(_1149_),
    .B(_0439_),
    .Y(_2792_));
 INVx2_ASAP7_75t_R _6042_ (.A(_2792_),
    .Y(_3136_));
 INVx2_ASAP7_75t_R _6043_ (.A(_1355_),
    .Y(_3157_));
 INVx2_ASAP7_75t_R _6044_ (.A(_3463_),
    .Y(_3464_));
 INVx2_ASAP7_75t_R _6045_ (.A(_1375_),
    .Y(_3160_));
 INVx2_ASAP7_75t_R _6046_ (.A(_3472_),
    .Y(_3473_));
 INVx2_ASAP7_75t_R _6047_ (.A(_1402_),
    .Y(_3163_));
 OR3x2_ASAP7_75t_R _6048_ (.A(_0352_),
    .B(_0366_),
    .C(_2768_),
    .Y(_2793_));
 OA21x2_ASAP7_75t_R _6049_ (.A1(_0356_),
    .A2(_0352_),
    .B(_0350_),
    .Y(_2794_));
 NAND2x2_ASAP7_75t_R _6050_ (.A(_2793_),
    .B(_2794_),
    .Y(_3140_));
 NAND2x2_ASAP7_75t_R _6051_ (.A(_0389_),
    .B(_2765_),
    .Y(_3144_));
 OA21x2_ASAP7_75t_R _6052_ (.A1(_0476_),
    .A2(_1524_),
    .B(_0001_),
    .Y(_2795_));
 OA21x2_ASAP7_75t_R _6053_ (.A1(net165),
    .A2(_2795_),
    .B(_0000_),
    .Y(_2796_));
 INVx2_ASAP7_75t_R _6054_ (.A(_2796_),
    .Y(_3153_));
 INVx2_ASAP7_75t_R _6055_ (.A(_1524_),
    .Y(_3158_));
 INVx2_ASAP7_75t_R _6056_ (.A(_1522_),
    .Y(_3161_));
 INVx2_ASAP7_75t_R _6057_ (.A(_1573_),
    .Y(_3522_));
 INVx2_ASAP7_75t_R _6058_ (.A(_1520_),
    .Y(_3164_));
 INVx2_ASAP7_75t_R _6059_ (.A(_1578_),
    .Y(_3527_));
 OA21x2_ASAP7_75t_R _6060_ (.A1(_0467_),
    .A2(_1518_),
    .B(_0009_),
    .Y(_2797_));
 OA21x2_ASAP7_75t_R _6061_ (.A1(net185),
    .A2(_2797_),
    .B(_0008_),
    .Y(_2798_));
 INVx2_ASAP7_75t_R _6062_ (.A(_2798_),
    .Y(_3167_));
 INVx2_ASAP7_75t_R _6063_ (.A(_1583_),
    .Y(_3532_));
 INVx2_ASAP7_75t_R _6064_ (.A(_1518_),
    .Y(_3170_));
 INVx2_ASAP7_75t_R _6065_ (.A(_1588_),
    .Y(_3537_));
 INVx2_ASAP7_75t_R _6066_ (.A(_1590_),
    .Y(_3181_));
 INVx2_ASAP7_75t_R _6067_ (.A(_1592_),
    .Y(_3177_));
 OR2x2_ASAP7_75t_R _6068_ (.A(_1594_),
    .B(_1677_),
    .Y(_2799_));
 OA21x2_ASAP7_75t_R _6069_ (.A1(_0748_),
    .A2(net221),
    .B(_2799_),
    .Y(_3545_));
 OA21x2_ASAP7_75t_R _6070_ (.A1(_0047_),
    .A2(_1697_),
    .B(_0065_),
    .Y(_2800_));
 OA21x2_ASAP7_75t_R _6071_ (.A1(net231),
    .A2(_2800_),
    .B(_0064_),
    .Y(_2801_));
 INVx2_ASAP7_75t_R _6072_ (.A(_2801_),
    .Y(_3184_));
 AND2x2_ASAP7_75t_R _6073_ (.A(_1580_),
    .B(net225),
    .Y(_2802_));
 AO21x2_ASAP7_75t_R _6074_ (.A1(_0068_),
    .A2(_1677_),
    .B(_2802_),
    .Y(_3550_));
 INVx2_ASAP7_75t_R _6075_ (.A(_1697_),
    .Y(_3187_));
 AND2x2_ASAP7_75t_R _6076_ (.A(_1585_),
    .B(net225),
    .Y(_2803_));
 AO21x2_ASAP7_75t_R _6077_ (.A1(_0071_),
    .A2(_1677_),
    .B(_2803_),
    .Y(_3552_));
 AND2x2_ASAP7_75t_R _6078_ (.A(_1564_),
    .B(net221),
    .Y(_2804_));
 AO21x2_ASAP7_75t_R _6079_ (.A1(_0082_),
    .A2(_1677_),
    .B(_2804_),
    .Y(_3555_));
 XOR2x2_ASAP7_75t_R _6080_ (.A(_0742_),
    .B(_0573_),
    .Y(_2805_));
 OR2x2_ASAP7_75t_R _6081_ (.A(_1676_),
    .B(_2805_),
    .Y(_2806_));
 OA21x2_ASAP7_75t_R _6082_ (.A1(_1568_),
    .A2(_1677_),
    .B(_2806_),
    .Y(_3556_));
 AND2x2_ASAP7_75t_R _6083_ (.A(_1570_),
    .B(_1676_),
    .Y(_2807_));
 AO21x2_ASAP7_75t_R _6084_ (.A1(_0574_),
    .A2(_1677_),
    .B(_2807_),
    .Y(_3557_));
 INVx2_ASAP7_75t_R _6085_ (.A(_1699_),
    .Y(_3196_));
 AND2x2_ASAP7_75t_R _6086_ (.A(_1575_),
    .B(_1676_),
    .Y(_2808_));
 AO21x2_ASAP7_75t_R _6087_ (.A1(_0086_),
    .A2(_1677_),
    .B(_2808_),
    .Y(_3559_));
 INVx2_ASAP7_75t_R _6088_ (.A(_1870_),
    .Y(_3581_));
 NOR2x2_ASAP7_75t_R _6089_ (.A(_1879_),
    .B(_1883_),
    .Y(_3583_));
 OR2x2_ASAP7_75t_R _6090_ (.A(_0119_),
    .B(net228),
    .Y(_2809_));
 NAND2x2_ASAP7_75t_R _6091_ (.A(_2809_),
    .B(_1884_),
    .Y(_3585_));
 INVx2_ASAP7_75t_R _6092_ (.A(_1921_),
    .Y(_3600_));
 NOR2x2_ASAP7_75t_R _6093_ (.A(_1916_),
    .B(_1918_),
    .Y(_3222_));
 AO21x2_ASAP7_75t_R _6094_ (.A1(_1927_),
    .A2(_1855_),
    .B(_1893_),
    .Y(_2810_));
 OA21x2_ASAP7_75t_R _6095_ (.A1(net219),
    .A2(_2005_),
    .B(_2810_),
    .Y(_2811_));
 OA21x2_ASAP7_75t_R _6096_ (.A1(_0162_),
    .A2(_3237_),
    .B(_0161_),
    .Y(_2812_));
 NOR2x2_ASAP7_75t_R _6097_ (.A(_2811_),
    .B(_2812_),
    .Y(_3612_));
 OA211x2_ASAP7_75t_R _6098_ (.A1(_2067_),
    .A2(_2068_),
    .B(_3612_),
    .C(_3611_),
    .Y(_3610_));
 INVx2_ASAP7_75t_R _6099_ (.A(_1965_),
    .Y(_3241_));
 INVx2_ASAP7_75t_R _6100_ (.A(_1940_),
    .Y(_3246_));
 AND4x2_ASAP7_75t_R _6101_ (.A(_2065_),
    .B(_2069_),
    .C(_3619_),
    .D(_2055_),
    .Y(_3615_));
 AO21x2_ASAP7_75t_R _6102_ (.A1(_0202_),
    .A2(_2155_),
    .B(_0201_),
    .Y(_2813_));
 NAND2x2_ASAP7_75t_R _6103_ (.A(_0794_),
    .B(_2813_),
    .Y(_3261_));
 AND2x2_ASAP7_75t_R _6104_ (.A(_2148_),
    .B(_2149_),
    .Y(_2814_));
 NOR2x2_ASAP7_75t_R _6105_ (.A(_2814_),
    .B(_2151_),
    .Y(_3264_));
 OR2x2_ASAP7_75t_R _6106_ (.A(_0799_),
    .B(_2144_),
    .Y(_2815_));
 OA21x2_ASAP7_75t_R _6107_ (.A1(_2142_),
    .A2(_2815_),
    .B(_0216_),
    .Y(_2816_));
 INVx2_ASAP7_75t_R _6108_ (.A(_2816_),
    .Y(_3284_));
 INVx2_ASAP7_75t_R _6109_ (.A(_2171_),
    .Y(_3649_));
 INVx2_ASAP7_75t_R _6110_ (.A(_2504_),
    .Y(_3306_));
 INVx2_ASAP7_75t_R _6111_ (.A(_2718_),
    .Y(_3671_));
 INVx2_ASAP7_75t_R _6112_ (.A(_2524_),
    .Y(_3319_));
 OA21x2_ASAP7_75t_R _6113_ (.A1(_0833_),
    .A2(_2520_),
    .B(_0295_),
    .Y(_2817_));
 INVx2_ASAP7_75t_R _6114_ (.A(_2817_),
    .Y(_3322_));
 INVx2_ASAP7_75t_R _6115_ (.A(_2519_),
    .Y(_3324_));
 INVx2_ASAP7_75t_R _6116_ (.A(_2560_),
    .Y(_3346_));
 INVx2_ASAP7_75t_R _6117_ (.A(_2517_),
    .Y(_3327_));
 INVx2_ASAP7_75t_R _6118_ (.A(_2532_),
    .Y(_3678_));
 OA21x2_ASAP7_75t_R _6119_ (.A1(_0309_),
    .A2(_3336_),
    .B(_0308_),
    .Y(_2818_));
 NOR2x2_ASAP7_75t_R _6120_ (.A(_2643_),
    .B(_2818_),
    .Y(_3681_));
 INVx2_ASAP7_75t_R _6121_ (.A(_2540_),
    .Y(_3341_));
 INVx2_ASAP7_75t_R _6122_ (.A(_2538_),
    .Y(_3344_));
 INVx2_ASAP7_75t_R _6123_ (.A(_2536_),
    .Y(_3347_));
 INVx2_ASAP7_75t_R _6124_ (.A(_2534_),
    .Y(_3350_));
 OA21x2_ASAP7_75t_R _6125_ (.A1(_2576_),
    .A2(net221),
    .B(_2579_),
    .Y(_3682_));
 AND2x2_ASAP7_75t_R _6126_ (.A(_0663_),
    .B(_1877_),
    .Y(_2819_));
 AND2x2_ASAP7_75t_R _6127_ (.A(_0849_),
    .B(net180),
    .Y(_2820_));
 XNOR2x2_ASAP7_75t_R _6128_ (.A(_2643_),
    .B(_2820_),
    .Y(_2821_));
 XNOR2x2_ASAP7_75t_R _6129_ (.A(_2819_),
    .B(_2821_),
    .Y(_3687_));
 AO21x2_ASAP7_75t_R _6130_ (.A1(_1877_),
    .A2(_2629_),
    .B(_2668_),
    .Y(_2822_));
 AND2x2_ASAP7_75t_R _6131_ (.A(_3701_),
    .B(_2822_),
    .Y(_3697_));
 NAND2x2_ASAP7_75t_R _6132_ (.A(_2653_),
    .B(_2657_),
    .Y(_2823_));
 AND3x2_ASAP7_75t_R _6133_ (.A(_3680_),
    .B(_2823_),
    .C(_3681_),
    .Y(_3714_));
 CKINVDCx8_ASAP7_75t_R _6134_ (.A(_3357_),
    .Y(_3365_));
 AND2x2_ASAP7_75t_R _6135_ (.A(_3685_),
    .B(_2726_),
    .Y(_3717_));
 OA211x2_ASAP7_75t_R _6136_ (.A1(_2740_),
    .A2(_2741_),
    .B(_2743_),
    .C(_0395_),
    .Y(_2824_));
 INVx2_ASAP7_75t_R _6137_ (.A(_2824_),
    .Y(_3366_));
 AND2x2_ASAP7_75t_R _6138_ (.A(_2715_),
    .B(_2735_),
    .Y(_2825_));
 NOR2x2_ASAP7_75t_R _6139_ (.A(_2825_),
    .B(_2733_),
    .Y(_3372_));
 INVx2_ASAP7_75t_R _6140_ (.A(_0427_),
    .Y(_2826_));
 NAND2x2_ASAP7_75t_R _6141_ (.A(_2826_),
    .B(_2754_),
    .Y(_2827_));
 TAPCELL_ASAP7_75t_R PHY_48 ();
 AND2x2_ASAP7_75t_R _6143_ (.A(\__st_1[0] ),
    .B(_2827_),
    .Y(_2829_));
 NAND3x2_ASAP7_75t_R _6144_ (.B(_2069_),
    .C(_2055_),
    .Y(_2830_),
    .A(_2065_));
 AND2x6_ASAP7_75t_R _6145_ (.A(_2826_),
    .B(_2754_),
    .Y(_2831_));
 XNOR2x2_ASAP7_75t_R _6146_ (.A(_0567_),
    .B(_0610_),
    .Y(_2832_));
 NOR2x2_ASAP7_75t_R _6147_ (.A(net162),
    .B(_2832_),
    .Y(_2833_));
 OA211x2_ASAP7_75t_R _6148_ (.A1(_2053_),
    .A2(_2830_),
    .B(_2831_),
    .C(_2833_),
    .Y(_2834_));
 AND4x2_ASAP7_75t_R _6149_ (.A(_2055_),
    .B(_2071_),
    .C(_2831_),
    .D(_2832_),
    .Y(_2835_));
 OA21x2_ASAP7_75t_R _6150_ (.A1(_1857_),
    .A2(_1863_),
    .B(_3609_),
    .Y(_2836_));
 INVx2_ASAP7_75t_R _6151_ (.A(_0180_),
    .Y(_2837_));
 OA211x2_ASAP7_75t_R _6152_ (.A1(_2074_),
    .A2(_2837_),
    .B(_1956_),
    .C(_1961_),
    .Y(_2838_));
 OA21x2_ASAP7_75t_R _6153_ (.A1(_2836_),
    .A2(_2838_),
    .B(_2833_),
    .Y(_2839_));
 AND2x2_ASAP7_75t_R _6154_ (.A(net162),
    .B(_2832_),
    .Y(_2840_));
 OA21x2_ASAP7_75t_R _6155_ (.A1(_2839_),
    .A2(_2840_),
    .B(_2831_),
    .Y(_2841_));
 AO21x2_ASAP7_75t_R _6156_ (.A1(_3619_),
    .A2(_2835_),
    .B(_2841_),
    .Y(_2842_));
 OR2x6_ASAP7_75t_R _6157_ (.A(_2834_),
    .B(_2842_),
    .Y(_2843_));
 TAPCELL_ASAP7_75t_R PHY_47 ();
 TAPCELL_ASAP7_75t_R PHY_46 ();
 INVx2_ASAP7_75t_R _6160_ (.A(_0242_),
    .Y(_2846_));
 AND4x2_ASAP7_75t_R _6161_ (.A(_2846_),
    .B(_0621_),
    .C(_0619_),
    .D(_0611_),
    .Y(_2847_));
 AND4x2_ASAP7_75t_R _6162_ (.A(_0617_),
    .B(_0623_),
    .C(_0615_),
    .D(_0613_),
    .Y(_2848_));
 XOR2x2_ASAP7_75t_R _6163_ (.A(_0189_),
    .B(_0612_),
    .Y(_2849_));
 XOR2x2_ASAP7_75t_R _6164_ (.A(_0241_),
    .B(_0796_),
    .Y(_2850_));
 XNOR2x2_ASAP7_75t_R _6165_ (.A(_0795_),
    .B(_0622_),
    .Y(_2851_));
 XNOR2x2_ASAP7_75t_R _6166_ (.A(_0618_),
    .B(_0793_),
    .Y(_2852_));
 AND4x2_ASAP7_75t_R _6167_ (.A(_2849_),
    .B(_2850_),
    .C(_2851_),
    .D(_2852_),
    .Y(_2853_));
 XNOR2x2_ASAP7_75t_R _6168_ (.A(_0798_),
    .B(_0637_),
    .Y(_2854_));
 XOR2x2_ASAP7_75t_R _6169_ (.A(_0201_),
    .B(_0620_),
    .Y(_2855_));
 XOR2x2_ASAP7_75t_R _6170_ (.A(_0192_),
    .B(_0614_),
    .Y(_2856_));
 XOR2x2_ASAP7_75t_R _6171_ (.A(_0195_),
    .B(_0616_),
    .Y(_2857_));
 AND4x2_ASAP7_75t_R _6172_ (.A(_2854_),
    .B(_2855_),
    .C(_2856_),
    .D(_2857_),
    .Y(_2858_));
 AND4x2_ASAP7_75t_R _6173_ (.A(_2847_),
    .B(_2848_),
    .C(_2853_),
    .D(_2858_),
    .Y(_2859_));
 INVx2_ASAP7_75t_R _6174_ (.A(_2859_),
    .Y(_2860_));
 OA211x2_ASAP7_75t_R _6175_ (.A1(_2053_),
    .A2(_2072_),
    .B(_2833_),
    .C(_2860_),
    .Y(_2861_));
 TAPCELL_ASAP7_75t_R PHY_45 ();
 AND4x2_ASAP7_75t_R _6177_ (.A(_2055_),
    .B(_2071_),
    .C(_2832_),
    .D(_2860_),
    .Y(_2863_));
 AO22x2_ASAP7_75t_R _6178_ (.A1(_2840_),
    .A2(_2860_),
    .B1(_2863_),
    .B2(_3619_),
    .Y(_2864_));
 TAPCELL_ASAP7_75t_R PHY_44 ();
 OR3x2_ASAP7_75t_R _6180_ (.A(_2855_),
    .B(_2851_),
    .C(_2856_),
    .Y(_2866_));
 OR4x2_ASAP7_75t_R _6181_ (.A(_0621_),
    .B(_0619_),
    .C(_0617_),
    .D(_0611_),
    .Y(_2867_));
 OR5x2_ASAP7_75t_R _6182_ (.A(_2846_),
    .B(_0623_),
    .C(_0615_),
    .D(_0613_),
    .E(_2867_),
    .Y(_2868_));
 OR4x2_ASAP7_75t_R _6183_ (.A(_2854_),
    .B(_2850_),
    .C(_2852_),
    .D(_2857_),
    .Y(_2869_));
 OR5x2_ASAP7_75t_R _6184_ (.A(_2827_),
    .B(_2849_),
    .C(_2866_),
    .D(_2868_),
    .E(_2869_),
    .Y(_2870_));
 NOR3x2_ASAP7_75t_R _6185_ (.B(_2864_),
    .C(_2870_),
    .Y(_2871_),
    .A(_2861_));
 TAPCELL_ASAP7_75t_R PHY_43 ();
 TAPCELL_ASAP7_75t_R PHY_42 ();
 TAPCELL_ASAP7_75t_R PHY_41 ();
 OR2x2_ASAP7_75t_R _6189_ (.A(_0120_),
    .B(_2829_),
    .Y(_2875_));
 CKINVDCx20_ASAP7_75t_R _6190_ (.A(net19),
    .Y(_2876_));
 TAPCELL_ASAP7_75t_R PHY_40 ();
 OA31x2_ASAP7_75t_R _6192_ (.A1(_2861_),
    .A2(_2864_),
    .A3(_2875_),
    .B1(_2876_),
    .Y(_2878_));
 OA31x2_ASAP7_75t_R _6193_ (.A1(_2829_),
    .A2(_2843_),
    .A3(net224),
    .B1(_2878_),
    .Y(_0869_));
 INVx2_ASAP7_75t_R _6194_ (.A(_3123_),
    .Y(_2879_));
 AND2x2_ASAP7_75t_R _6195_ (.A(_2879_),
    .B(_2827_),
    .Y(_2880_));
 OR2x2_ASAP7_75t_R _6196_ (.A(_0624_),
    .B(_2880_),
    .Y(_2881_));
 OA31x2_ASAP7_75t_R _6197_ (.A1(_2861_),
    .A2(_2864_),
    .A3(_2881_),
    .B1(_2876_),
    .Y(_2882_));
 OA31x2_ASAP7_75t_R _6198_ (.A1(_2843_),
    .A2(net224),
    .A3(_2880_),
    .B1(_2882_),
    .Y(_0870_));
 AND2x2_ASAP7_75t_R _6199_ (.A(\__st_1[2] ),
    .B(_2827_),
    .Y(_2883_));
 OR2x2_ASAP7_75t_R _6200_ (.A(_0626_),
    .B(_2883_),
    .Y(_2884_));
 OA31x2_ASAP7_75t_R _6201_ (.A1(_2861_),
    .A2(_2864_),
    .A3(_2884_),
    .B1(_2876_),
    .Y(_2885_));
 OA31x2_ASAP7_75t_R _6202_ (.A1(_2843_),
    .A2(net224),
    .A3(_2883_),
    .B1(_2885_),
    .Y(_0871_));
 TAPCELL_ASAP7_75t_R PHY_39 ();
 AND2x2_ASAP7_75t_R _6204_ (.A(\__st_1[3] ),
    .B(_2827_),
    .Y(_2887_));
 XNOR2x2_ASAP7_75t_R _6205_ (.A(_0625_),
    .B(_0809_),
    .Y(_2888_));
 OR2x2_ASAP7_75t_R _6206_ (.A(_2887_),
    .B(_2888_),
    .Y(_2889_));
 OA31x2_ASAP7_75t_R _6207_ (.A1(_2861_),
    .A2(_2864_),
    .A3(_2889_),
    .B1(_2876_),
    .Y(_2890_));
 OA31x2_ASAP7_75t_R _6208_ (.A1(_2843_),
    .A2(net224),
    .A3(_2887_),
    .B1(_2890_),
    .Y(_0872_));
 AND2x2_ASAP7_75t_R _6209_ (.A(\__st_1[4] ),
    .B(_2827_),
    .Y(_2891_));
 OR2x2_ASAP7_75t_R _6210_ (.A(_0628_),
    .B(_2891_),
    .Y(_2892_));
 TAPCELL_ASAP7_75t_R PHY_38 ();
 OA31x2_ASAP7_75t_R _6212_ (.A1(_2861_),
    .A2(_2864_),
    .A3(_2892_),
    .B1(_2876_),
    .Y(_2894_));
 OA31x2_ASAP7_75t_R _6213_ (.A1(_2843_),
    .A2(net224),
    .A3(_2891_),
    .B1(_2894_),
    .Y(_0873_));
 AND2x2_ASAP7_75t_R _6214_ (.A(\__st_1[5] ),
    .B(_2827_),
    .Y(_2895_));
 XNOR2x2_ASAP7_75t_R _6215_ (.A(_0807_),
    .B(_0627_),
    .Y(_2896_));
 OR2x2_ASAP7_75t_R _6216_ (.A(_2895_),
    .B(_2896_),
    .Y(_2897_));
 OA31x2_ASAP7_75t_R _6217_ (.A1(_2861_),
    .A2(_2864_),
    .A3(_2897_),
    .B1(_2876_),
    .Y(_2898_));
 OA31x2_ASAP7_75t_R _6218_ (.A1(_2843_),
    .A2(net235),
    .A3(_2895_),
    .B1(_2898_),
    .Y(_0874_));
 AND2x2_ASAP7_75t_R _6219_ (.A(\__st_1[6] ),
    .B(_2827_),
    .Y(_2899_));
 OR2x2_ASAP7_75t_R _6220_ (.A(_0630_),
    .B(_2899_),
    .Y(_2900_));
 OA31x2_ASAP7_75t_R _6221_ (.A1(_2861_),
    .A2(_2864_),
    .A3(_2900_),
    .B1(_2876_),
    .Y(_2901_));
 OA31x2_ASAP7_75t_R _6222_ (.A1(_2843_),
    .A2(net235),
    .A3(_2899_),
    .B1(_2901_),
    .Y(_0875_));
 AND2x2_ASAP7_75t_R _6223_ (.A(\__st_1[7] ),
    .B(_2827_),
    .Y(_2902_));
 XNOR2x2_ASAP7_75t_R _6224_ (.A(_0805_),
    .B(_0629_),
    .Y(_2903_));
 OR2x2_ASAP7_75t_R _6225_ (.A(_2902_),
    .B(_2903_),
    .Y(_2904_));
 OA31x2_ASAP7_75t_R _6226_ (.A1(_2861_),
    .A2(_2864_),
    .A3(_2904_),
    .B1(_2876_),
    .Y(_2905_));
 OA31x2_ASAP7_75t_R _6227_ (.A1(_2843_),
    .A2(net235),
    .A3(_2902_),
    .B1(_2905_),
    .Y(_0876_));
 AND2x2_ASAP7_75t_R _6228_ (.A(\__st_1[8] ),
    .B(_2827_),
    .Y(_2906_));
 OR2x2_ASAP7_75t_R _6229_ (.A(_0632_),
    .B(_2906_),
    .Y(_2907_));
 OA31x2_ASAP7_75t_R _6230_ (.A1(_2861_),
    .A2(_2864_),
    .A3(_2907_),
    .B1(_2876_),
    .Y(_2908_));
 OA31x2_ASAP7_75t_R _6231_ (.A1(_2843_),
    .A2(net235),
    .A3(_2906_),
    .B1(_2908_),
    .Y(_0877_));
 AND2x2_ASAP7_75t_R _6232_ (.A(\__st_1[9] ),
    .B(_2827_),
    .Y(_2909_));
 XNOR2x2_ASAP7_75t_R _6233_ (.A(_0803_),
    .B(_0631_),
    .Y(_2910_));
 OR2x2_ASAP7_75t_R _6234_ (.A(_2909_),
    .B(_2910_),
    .Y(_2911_));
 OA31x2_ASAP7_75t_R _6235_ (.A1(_2861_),
    .A2(_2864_),
    .A3(_2911_),
    .B1(_2876_),
    .Y(_2912_));
 OA31x2_ASAP7_75t_R _6236_ (.A1(_2843_),
    .A2(net235),
    .A3(_2909_),
    .B1(_2912_),
    .Y(_0878_));
 AND2x2_ASAP7_75t_R _6237_ (.A(\__st_1[10] ),
    .B(_2827_),
    .Y(_2913_));
 OR2x2_ASAP7_75t_R _6238_ (.A(_0634_),
    .B(_2913_),
    .Y(_2914_));
 OA31x2_ASAP7_75t_R _6239_ (.A1(_2861_),
    .A2(_2864_),
    .A3(_2914_),
    .B1(_2876_),
    .Y(_2915_));
 OA31x2_ASAP7_75t_R _6240_ (.A1(_2843_),
    .A2(net235),
    .A3(_2913_),
    .B1(_2915_),
    .Y(_0879_));
 AND2x2_ASAP7_75t_R _6241_ (.A(\__st_1[11] ),
    .B(_2827_),
    .Y(_2916_));
 XNOR2x2_ASAP7_75t_R _6242_ (.A(_0801_),
    .B(_0633_),
    .Y(_2917_));
 OR2x2_ASAP7_75t_R _6243_ (.A(_2916_),
    .B(_2917_),
    .Y(_2918_));
 OA31x2_ASAP7_75t_R _6244_ (.A1(_2861_),
    .A2(_2864_),
    .A3(_2918_),
    .B1(_2876_),
    .Y(_2919_));
 OA31x2_ASAP7_75t_R _6245_ (.A1(_2843_),
    .A2(net235),
    .A3(_2916_),
    .B1(_2919_),
    .Y(_0880_));
 AND2x2_ASAP7_75t_R _6246_ (.A(\__st_1[12] ),
    .B(_2827_),
    .Y(_2920_));
 OR2x2_ASAP7_75t_R _6247_ (.A(_0636_),
    .B(_2920_),
    .Y(_2921_));
 OA31x2_ASAP7_75t_R _6248_ (.A1(_2861_),
    .A2(_2864_),
    .A3(_2921_),
    .B1(_2876_),
    .Y(_2922_));
 OA31x2_ASAP7_75t_R _6249_ (.A1(_2843_),
    .A2(net235),
    .A3(_2920_),
    .B1(_2922_),
    .Y(_0881_));
 AND2x2_ASAP7_75t_R _6250_ (.A(\__st_1[13] ),
    .B(_2827_),
    .Y(_2923_));
 XNOR2x2_ASAP7_75t_R _6251_ (.A(_0799_),
    .B(_0635_),
    .Y(_2924_));
 OR2x2_ASAP7_75t_R _6252_ (.A(_2923_),
    .B(_2924_),
    .Y(_2925_));
 OA31x2_ASAP7_75t_R _6253_ (.A1(_2861_),
    .A2(_2864_),
    .A3(_2925_),
    .B1(_2876_),
    .Y(_2926_));
 OA31x2_ASAP7_75t_R _6254_ (.A1(_2843_),
    .A2(net224),
    .A3(_2923_),
    .B1(_2926_),
    .Y(_0882_));
 AND2x2_ASAP7_75t_R _6255_ (.A(\__st_1[14] ),
    .B(_2827_),
    .Y(_2927_));
 OR2x2_ASAP7_75t_R _6256_ (.A(_0638_),
    .B(_2927_),
    .Y(_2928_));
 OA31x2_ASAP7_75t_R _6257_ (.A1(_2861_),
    .A2(_2864_),
    .A3(_2928_),
    .B1(_2876_),
    .Y(_2929_));
 OA31x2_ASAP7_75t_R _6258_ (.A1(_2843_),
    .A2(net224),
    .A3(_2927_),
    .B1(_2929_),
    .Y(_0883_));
 TAPCELL_ASAP7_75t_R PHY_37 ();
 TAPCELL_ASAP7_75t_R PHY_36 ();
 TAPCELL_ASAP7_75t_R PHY_35 ();
 NOR3x2_ASAP7_75t_R _6262_ (.B(_2834_),
    .C(_2842_),
    .Y(_2933_),
    .A(net19));
 TAPCELL_ASAP7_75t_R PHY_34 ();
 OA21x2_ASAP7_75t_R _6264_ (.A1(\__st_1[15] ),
    .A2(_2831_),
    .B(_2933_),
    .Y(_0884_));
 OA21x2_ASAP7_75t_R _6265_ (.A1(\__st_1[16] ),
    .A2(_2831_),
    .B(_2933_),
    .Y(_0885_));
 OA21x2_ASAP7_75t_R _6266_ (.A1(\__st_1[17] ),
    .A2(_2831_),
    .B(_2933_),
    .Y(_0886_));
 OA21x2_ASAP7_75t_R _6267_ (.A1(\__st_1[18] ),
    .A2(_2831_),
    .B(_2933_),
    .Y(_0887_));
 OA21x2_ASAP7_75t_R _6268_ (.A1(\__st_1[19] ),
    .A2(_2831_),
    .B(_2933_),
    .Y(_0888_));
 OA21x2_ASAP7_75t_R _6269_ (.A1(\__st_1[20] ),
    .A2(_2831_),
    .B(_2933_),
    .Y(_0889_));
 OA21x2_ASAP7_75t_R _6270_ (.A1(\__st_1[21] ),
    .A2(_2831_),
    .B(_2933_),
    .Y(_0890_));
 OA21x2_ASAP7_75t_R _6271_ (.A1(\__st_1[22] ),
    .A2(_2831_),
    .B(_2933_),
    .Y(_0891_));
 OA21x2_ASAP7_75t_R _6272_ (.A1(\__st_1[23] ),
    .A2(_2831_),
    .B(_2933_),
    .Y(_0892_));
 OA21x2_ASAP7_75t_R _6273_ (.A1(\__st_1[24] ),
    .A2(_2831_),
    .B(_2933_),
    .Y(_0893_));
 TAPCELL_ASAP7_75t_R PHY_33 ();
 TAPCELL_ASAP7_75t_R PHY_32 ();
 OA21x2_ASAP7_75t_R _6276_ (.A1(\__st_1[25] ),
    .A2(_2831_),
    .B(_2933_),
    .Y(_0894_));
 OA21x2_ASAP7_75t_R _6277_ (.A1(\__st_1[26] ),
    .A2(_2831_),
    .B(_2933_),
    .Y(_0895_));
 OA21x2_ASAP7_75t_R _6278_ (.A1(\__st_1[27] ),
    .A2(_2831_),
    .B(_2933_),
    .Y(_0896_));
 OA21x2_ASAP7_75t_R _6279_ (.A1(\__st_1[28] ),
    .A2(_2831_),
    .B(_2933_),
    .Y(_0897_));
 OA21x2_ASAP7_75t_R _6280_ (.A1(\__st_1[29] ),
    .A2(_2831_),
    .B(_2933_),
    .Y(_0898_));
 INVx2_ASAP7_75t_R _6281_ (.A(_3139_),
    .Y(_2937_));
 OA21x2_ASAP7_75t_R _6282_ (.A1(_2937_),
    .A2(_2831_),
    .B(_2933_),
    .Y(_0899_));
 OA21x2_ASAP7_75t_R _6283_ (.A1(_1171_),
    .A2(_2831_),
    .B(_2933_),
    .Y(_0900_));
 TAPCELL_ASAP7_75t_R PHY_31 ();
 TAPCELL_ASAP7_75t_R PHY_30 ();
 XNOR2x2_ASAP7_75t_R _6286_ (.A(_0639_),
    .B(net229),
    .Y(_2940_));
 INVx2_ASAP7_75t_R _6287_ (.A(_0648_),
    .Y(_2941_));
 AND3x2_ASAP7_75t_R _6288_ (.A(_0264_),
    .B(_2941_),
    .C(_0813_),
    .Y(_2942_));
 XOR2x2_ASAP7_75t_R _6289_ (.A(_0647_),
    .B(_0816_),
    .Y(_2943_));
 OR2x2_ASAP7_75t_R _6290_ (.A(_0262_),
    .B(_2943_),
    .Y(_2944_));
 XNOR2x2_ASAP7_75t_R _6291_ (.A(_0261_),
    .B(_0562_),
    .Y(_2945_));
 OA21x2_ASAP7_75t_R _6292_ (.A1(_2942_),
    .A2(_2944_),
    .B(_2945_),
    .Y(_2946_));
 XNOR2x2_ASAP7_75t_R _6293_ (.A(_0639_),
    .B(net38),
    .Y(_2947_));
 OR2x2_ASAP7_75t_R _6294_ (.A(_0260_),
    .B(_2947_),
    .Y(_2948_));
 XOR2x2_ASAP7_75t_R _6295_ (.A(_0255_),
    .B(_0817_),
    .Y(_2949_));
 OR5x2_ASAP7_75t_R _6296_ (.A(_0646_),
    .B(_0644_),
    .C(_0642_),
    .D(_0640_),
    .E(_2949_),
    .Y(_2950_));
 XNOR2x2_ASAP7_75t_R _6297_ (.A(_0641_),
    .B(_0814_),
    .Y(_2951_));
 XNOR2x2_ASAP7_75t_R _6298_ (.A(_0643_),
    .B(_0815_),
    .Y(_2952_));
 XOR2x2_ASAP7_75t_R _6299_ (.A(_0251_),
    .B(_0645_),
    .Y(_2953_));
 OR3x2_ASAP7_75t_R _6300_ (.A(_2951_),
    .B(_2952_),
    .C(_2953_),
    .Y(_2954_));
 OA21x2_ASAP7_75t_R _6301_ (.A1(_2950_),
    .A2(_2954_),
    .B(_2940_),
    .Y(_2955_));
 INVx2_ASAP7_75t_R _6302_ (.A(_2955_),
    .Y(_2956_));
 OA21x2_ASAP7_75t_R _6303_ (.A1(_2946_),
    .A2(_2948_),
    .B(_2956_),
    .Y(_2957_));
 AND2x2_ASAP7_75t_R _6304_ (.A(_2940_),
    .B(_2957_),
    .Y(_2958_));
 AND2x2_ASAP7_75t_R _6305_ (.A(_2831_),
    .B(_2958_),
    .Y(_2959_));
 INVx2_ASAP7_75t_R _6306_ (.A(_0813_),
    .Y(_2960_));
 AO22x2_ASAP7_75t_R _6307_ (.A1(\__st_2[0] ),
    .A2(_2827_),
    .B1(_2959_),
    .B2(_2960_),
    .Y(_2961_));
 AND2x2_ASAP7_75t_R _6308_ (.A(_2876_),
    .B(_2961_),
    .Y(_0901_));
 NAND2x2_ASAP7_75t_R _6309_ (.A(_2831_),
    .B(_2958_),
    .Y(_2962_));
 OA22x2_ASAP7_75t_R _6310_ (.A1(_0565_),
    .A2(_2831_),
    .B1(_2962_),
    .B2(_0264_),
    .Y(_2963_));
 NOR2x2_ASAP7_75t_R _6311_ (.A(net19),
    .B(_2963_),
    .Y(_0902_));
 AO22x2_ASAP7_75t_R _6312_ (.A1(\__st_2[2] ),
    .A2(_2827_),
    .B1(_2959_),
    .B2(_0648_),
    .Y(_2964_));
 AND2x2_ASAP7_75t_R _6313_ (.A(_2876_),
    .B(_2964_),
    .Y(_0903_));
 OA21x2_ASAP7_75t_R _6314_ (.A1(_2947_),
    .A2(_2943_),
    .B(_2957_),
    .Y(_2965_));
 AO21x2_ASAP7_75t_R _6315_ (.A1(_0564_),
    .A2(_2827_),
    .B(net19),
    .Y(_2966_));
 AO21x2_ASAP7_75t_R _6316_ (.A1(_2831_),
    .A2(_2965_),
    .B(_2966_),
    .Y(_2967_));
 INVx2_ASAP7_75t_R _6317_ (.A(_2967_),
    .Y(_0904_));
 TAPCELL_ASAP7_75t_R PHY_29 ();
 TAPCELL_ASAP7_75t_R PHY_28 ();
 OA21x2_ASAP7_75t_R _6320_ (.A1(_0262_),
    .A2(_2947_),
    .B(_2831_),
    .Y(_2970_));
 AO221x2_ASAP7_75t_R _6321_ (.A1(_0563_),
    .A2(_2827_),
    .B1(_2957_),
    .B2(_2970_),
    .C(net19),
    .Y(_2971_));
 INVx2_ASAP7_75t_R _6322_ (.A(_2971_),
    .Y(_0905_));
 AO21x2_ASAP7_75t_R _6323_ (.A1(_0261_),
    .A2(_2958_),
    .B(_2827_),
    .Y(_2972_));
 AND2x2_ASAP7_75t_R _6324_ (.A(_2189_),
    .B(_2972_),
    .Y(_2973_));
 INVx2_ASAP7_75t_R _6325_ (.A(_0261_),
    .Y(_2974_));
 AND3x2_ASAP7_75t_R _6326_ (.A(_2974_),
    .B(_0562_),
    .C(_2959_),
    .Y(_2975_));
 TAPCELL_ASAP7_75t_R PHY_27 ();
 OA21x2_ASAP7_75t_R _6328_ (.A1(_2973_),
    .A2(_2975_),
    .B(_2876_),
    .Y(_0906_));
 AND3x2_ASAP7_75t_R _6329_ (.A(_2831_),
    .B(_2956_),
    .C(_2948_),
    .Y(_2977_));
 AO21x2_ASAP7_75t_R _6330_ (.A1(_0259_),
    .A2(_2827_),
    .B(net19),
    .Y(_2978_));
 NOR2x2_ASAP7_75t_R _6331_ (.A(_2977_),
    .B(_2978_),
    .Y(_0907_));
 AND2x6_ASAP7_75t_R _6332_ (.A(_2876_),
    .B(_2827_),
    .Y(_2979_));
 TAPCELL_ASAP7_75t_R PHY_26 ();
 AND2x2_ASAP7_75t_R _6334_ (.A(\__st_2[7] ),
    .B(_2979_),
    .Y(_0908_));
 AND2x2_ASAP7_75t_R _6335_ (.A(\__st_2[8] ),
    .B(_2979_),
    .Y(_0909_));
 AND2x2_ASAP7_75t_R _6336_ (.A(\__st_2[9] ),
    .B(_2979_),
    .Y(_0910_));
 AND2x2_ASAP7_75t_R _6337_ (.A(\__st_2[10] ),
    .B(_2979_),
    .Y(_0911_));
 AND2x2_ASAP7_75t_R _6338_ (.A(\__st_2[11] ),
    .B(_2979_),
    .Y(_0912_));
 AND2x2_ASAP7_75t_R _6339_ (.A(\__st_2[12] ),
    .B(_2979_),
    .Y(_0913_));
 AND2x2_ASAP7_75t_R _6340_ (.A(\__st_2[13] ),
    .B(_2979_),
    .Y(_0914_));
 INVx2_ASAP7_75t_R _6341_ (.A(_3285_),
    .Y(_2981_));
 AND2x2_ASAP7_75t_R _6342_ (.A(_2981_),
    .B(_2979_),
    .Y(_0915_));
 XNOR2x2_ASAP7_75t_R _6343_ (.A(_0575_),
    .B(net229),
    .Y(_2982_));
 INVx2_ASAP7_75t_R _6344_ (.A(_2982_),
    .Y(_2983_));
 INVx2_ASAP7_75t_R _6345_ (.A(_0113_),
    .Y(_2984_));
 INVx2_ASAP7_75t_R _6346_ (.A(_0115_),
    .Y(_2985_));
 INVx2_ASAP7_75t_R _6347_ (.A(_0116_),
    .Y(_2986_));
 INVx2_ASAP7_75t_R _6348_ (.A(_0730_),
    .Y(_2987_));
 OR3x2_ASAP7_75t_R _6349_ (.A(_2986_),
    .B(_0584_),
    .C(_2987_),
    .Y(_2988_));
 XNOR2x2_ASAP7_75t_R _6350_ (.A(_0583_),
    .B(_0765_),
    .Y(_2989_));
 AND3x2_ASAP7_75t_R _6351_ (.A(_2985_),
    .B(_2988_),
    .C(_2989_),
    .Y(_2990_));
 XOR2x2_ASAP7_75t_R _6352_ (.A(_0114_),
    .B(_0552_),
    .Y(_2991_));
 AO21x2_ASAP7_75t_R _6353_ (.A1(_2982_),
    .A2(_2990_),
    .B(_2991_),
    .Y(_2992_));
 XOR2x2_ASAP7_75t_R _6354_ (.A(_0514_),
    .B(_0766_),
    .Y(_2993_));
 OR4x2_ASAP7_75t_R _6355_ (.A(_0580_),
    .B(_0578_),
    .C(_0576_),
    .D(_0582_),
    .Y(_2994_));
 XNOR2x2_ASAP7_75t_R _6356_ (.A(_0579_),
    .B(_0732_),
    .Y(_2995_));
 XNOR2x2_ASAP7_75t_R _6357_ (.A(_0577_),
    .B(_0731_),
    .Y(_2996_));
 XOR2x2_ASAP7_75t_R _6358_ (.A(_0510_),
    .B(_0581_),
    .Y(_2997_));
 OR5x2_ASAP7_75t_R _6359_ (.A(_2993_),
    .B(_2994_),
    .C(_2995_),
    .D(_2996_),
    .E(_2997_),
    .Y(_2998_));
 AO21x2_ASAP7_75t_R _6360_ (.A1(_2984_),
    .A2(_2992_),
    .B(_2998_),
    .Y(_2999_));
 OR3x4_ASAP7_75t_R _6361_ (.A(_2827_),
    .B(_2983_),
    .C(_2999_),
    .Y(_3000_));
 OA22x2_ASAP7_75t_R _6362_ (.A1(_0556_),
    .A2(_2831_),
    .B1(_3000_),
    .B2(_0730_),
    .Y(_3001_));
 NOR2x2_ASAP7_75t_R _6363_ (.A(net19),
    .B(_3001_),
    .Y(_0916_));
 OA22x2_ASAP7_75t_R _6364_ (.A1(_0555_),
    .A2(_2831_),
    .B1(_3000_),
    .B2(_0116_),
    .Y(_3002_));
 NOR2x2_ASAP7_75t_R _6365_ (.A(net19),
    .B(_3002_),
    .Y(_0917_));
 INVx2_ASAP7_75t_R _6366_ (.A(_0584_),
    .Y(_3003_));
 OA22x2_ASAP7_75t_R _6367_ (.A1(_3206_),
    .A2(_2831_),
    .B1(_3000_),
    .B2(_3003_),
    .Y(_3004_));
 NOR2x2_ASAP7_75t_R _6368_ (.A(net19),
    .B(_3004_),
    .Y(_0918_));
 TAPCELL_ASAP7_75t_R PHY_25 ();
 OA21x2_ASAP7_75t_R _6370_ (.A1(_2989_),
    .A2(_2999_),
    .B(_2982_),
    .Y(_3006_));
 OA21x2_ASAP7_75t_R _6371_ (.A1(\__st_0[3] ),
    .A2(_2831_),
    .B(_2876_),
    .Y(_3007_));
 OA21x2_ASAP7_75t_R _6372_ (.A1(_2827_),
    .A2(_3006_),
    .B(_3007_),
    .Y(_0919_));
 AND2x2_ASAP7_75t_R _6373_ (.A(\__st_0[4] ),
    .B(_2827_),
    .Y(_3008_));
 OA211x2_ASAP7_75t_R _6374_ (.A1(_2985_),
    .A2(_2999_),
    .B(_2982_),
    .C(_2831_),
    .Y(_3009_));
 OA21x2_ASAP7_75t_R _6375_ (.A1(_3008_),
    .A2(_3009_),
    .B(_2876_),
    .Y(_0920_));
 INVx2_ASAP7_75t_R _6376_ (.A(_0114_),
    .Y(_3010_));
 OA21x2_ASAP7_75t_R _6377_ (.A1(_3010_),
    .A2(_3000_),
    .B(_2831_),
    .Y(_3011_));
 OR3x2_ASAP7_75t_R _6378_ (.A(_0114_),
    .B(_1000_),
    .C(_3000_),
    .Y(_3012_));
 OA21x2_ASAP7_75t_R _6379_ (.A1(_0552_),
    .A2(_3011_),
    .B(_3012_),
    .Y(_3013_));
 NOR2x2_ASAP7_75t_R _6380_ (.A(net19),
    .B(_3013_),
    .Y(_0921_));
 AND2x2_ASAP7_75t_R _6381_ (.A(\__st_0[6] ),
    .B(_2827_),
    .Y(_3014_));
 OA211x2_ASAP7_75t_R _6382_ (.A1(_2984_),
    .A2(_2998_),
    .B(_2982_),
    .C(_2831_),
    .Y(_3015_));
 OA21x2_ASAP7_75t_R _6383_ (.A1(_3014_),
    .A2(_3015_),
    .B(_2876_),
    .Y(_0922_));
 AND2x2_ASAP7_75t_R _6384_ (.A(\__st_0[7] ),
    .B(_2979_),
    .Y(_0923_));
 AND2x2_ASAP7_75t_R _6385_ (.A(\__st_0[8] ),
    .B(_2979_),
    .Y(_0924_));
 TAPCELL_ASAP7_75t_R PHY_24 ();
 AND2x2_ASAP7_75t_R _6387_ (.A(\__st_0[9] ),
    .B(_2979_),
    .Y(_0925_));
 AND2x2_ASAP7_75t_R _6388_ (.A(\__st_0[10] ),
    .B(_2979_),
    .Y(_0926_));
 AND2x2_ASAP7_75t_R _6389_ (.A(\__st_0[11] ),
    .B(_2979_),
    .Y(_0927_));
 AND2x2_ASAP7_75t_R _6390_ (.A(\__st_0[12] ),
    .B(_2979_),
    .Y(_0928_));
 AND2x2_ASAP7_75t_R _6391_ (.A(\__st_0[13] ),
    .B(_2979_),
    .Y(_0929_));
 INVx2_ASAP7_75t_R _6392_ (.A(_3197_),
    .Y(_3017_));
 AND2x2_ASAP7_75t_R _6393_ (.A(_3017_),
    .B(_2979_),
    .Y(_0930_));
 XNOR2x2_ASAP7_75t_R _6394_ (.A(_0529_),
    .B(_0667_),
    .Y(_3018_));
 INVx2_ASAP7_75t_R _6395_ (.A(_0412_),
    .Y(_3019_));
 OR4x2_ASAP7_75t_R _6396_ (.A(_0676_),
    .B(_0674_),
    .C(_0672_),
    .D(_0670_),
    .Y(_3020_));
 OR5x2_ASAP7_75t_R _6397_ (.A(_3019_),
    .B(_0680_),
    .C(_0678_),
    .D(_0668_),
    .E(_3020_),
    .Y(_3021_));
 XOR2x2_ASAP7_75t_R _6398_ (.A(_0387_),
    .B(_0673_),
    .Y(_3022_));
 XOR2x2_ASAP7_75t_R _6399_ (.A(_0381_),
    .B(_0669_),
    .Y(_3023_));
 XNOR2x2_ASAP7_75t_R _6400_ (.A(_0403_),
    .B(_0411_),
    .Y(_3024_));
 XNOR2x2_ASAP7_75t_R _6401_ (.A(_0675_),
    .B(_0864_),
    .Y(_3025_));
 OR5x2_ASAP7_75t_R _6402_ (.A(_3021_),
    .B(_3022_),
    .C(_3023_),
    .D(_3024_),
    .E(_3025_),
    .Y(_3026_));
 XOR2x2_ASAP7_75t_R _6403_ (.A(_0679_),
    .B(_0866_),
    .Y(_3027_));
 XOR2x2_ASAP7_75t_R _6404_ (.A(_0344_),
    .B(_0694_),
    .Y(_3028_));
 XOR2x2_ASAP7_75t_R _6405_ (.A(_0677_),
    .B(_0865_),
    .Y(_3029_));
 XOR2x2_ASAP7_75t_R _6406_ (.A(_0384_),
    .B(_0671_),
    .Y(_3030_));
 OR4x2_ASAP7_75t_R _6407_ (.A(_3027_),
    .B(_3028_),
    .C(_3029_),
    .D(_3030_),
    .Y(_3031_));
 NOR2x2_ASAP7_75t_R _6408_ (.A(_3026_),
    .B(_3031_),
    .Y(_3032_));
 OR2x2_ASAP7_75t_R _6409_ (.A(_3018_),
    .B(_3032_),
    .Y(_3033_));
 XOR2x2_ASAP7_75t_R _6410_ (.A(_0529_),
    .B(_0667_),
    .Y(_3034_));
 OR4x2_ASAP7_75t_R _6411_ (.A(net162),
    .B(_2727_),
    .C(_3034_),
    .D(_3032_),
    .Y(_3035_));
 OA211x2_ASAP7_75t_R _6412_ (.A1(_3357_),
    .A2(_3033_),
    .B(_3035_),
    .C(_2831_),
    .Y(_3036_));
 TAPCELL_ASAP7_75t_R PHY_23 ();
 AND4x2_ASAP7_75t_R _6414_ (.A(_3019_),
    .B(_0680_),
    .C(_0678_),
    .D(_0668_),
    .Y(_3038_));
 AND4x2_ASAP7_75t_R _6415_ (.A(_0676_),
    .B(_0674_),
    .C(_0672_),
    .D(_0670_),
    .Y(_3039_));
 AND4x2_ASAP7_75t_R _6416_ (.A(_3022_),
    .B(_3023_),
    .C(_3024_),
    .D(_3025_),
    .Y(_3040_));
 AND4x2_ASAP7_75t_R _6417_ (.A(_3027_),
    .B(_3028_),
    .C(_3029_),
    .D(_3030_),
    .Y(_3041_));
 AND4x2_ASAP7_75t_R _6418_ (.A(_3038_),
    .B(_3039_),
    .C(_3040_),
    .D(_3041_),
    .Y(_3042_));
 OR2x2_ASAP7_75t_R _6419_ (.A(_3018_),
    .B(_3042_),
    .Y(_3043_));
 NOR3x2_ASAP7_75t_R _6420_ (.B(_2727_),
    .C(_3043_),
    .Y(_3044_),
    .A(net162));
 INVx2_ASAP7_75t_R _6421_ (.A(_3042_),
    .Y(_3045_));
 OA211x2_ASAP7_75t_R _6422_ (.A1(net162),
    .A2(_2727_),
    .B(_3018_),
    .C(_3045_),
    .Y(_3046_));
 TAPCELL_ASAP7_75t_R PHY_22 ();
 OR3x2_ASAP7_75t_R _6424_ (.A(_0414_),
    .B(_3044_),
    .C(_3046_),
    .Y(_3048_));
 AO32x2_ASAP7_75t_R _6425_ (.A1(_2876_),
    .A2(_3036_),
    .A3(_3048_),
    .B1(_2979_),
    .B2(net21),
    .Y(_0931_));
 OR3x2_ASAP7_75t_R _6426_ (.A(_0681_),
    .B(_3044_),
    .C(_3046_),
    .Y(_3049_));
 AO32x2_ASAP7_75t_R _6427_ (.A1(_2876_),
    .A2(_3036_),
    .A3(_3049_),
    .B1(_2979_),
    .B2(net28),
    .Y(_0932_));
 OA211x2_ASAP7_75t_R _6428_ (.A1(_3357_),
    .A2(_3033_),
    .B(_3035_),
    .C(_0683_),
    .Y(_3050_));
 OR3x2_ASAP7_75t_R _6429_ (.A(_2827_),
    .B(_3044_),
    .C(_3046_),
    .Y(_3051_));
 OA21x2_ASAP7_75t_R _6430_ (.A1(net29),
    .A2(_2831_),
    .B(_2876_),
    .Y(_3052_));
 OA21x2_ASAP7_75t_R _6431_ (.A1(_3050_),
    .A2(_3051_),
    .B(_3052_),
    .Y(_0933_));
 AND2x2_ASAP7_75t_R _6432_ (.A(net30),
    .B(_2827_),
    .Y(_3053_));
 XNOR2x2_ASAP7_75t_R _6433_ (.A(_0859_),
    .B(_0682_),
    .Y(_3054_));
 OR2x2_ASAP7_75t_R _6434_ (.A(_3053_),
    .B(_3054_),
    .Y(_3055_));
 OR2x6_ASAP7_75t_R _6435_ (.A(_3044_),
    .B(_3046_),
    .Y(_3056_));
 TAPCELL_ASAP7_75t_R PHY_21 ();
 OA221x2_ASAP7_75t_R _6437_ (.A1(_3036_),
    .A2(_3053_),
    .B1(_3055_),
    .B2(_3056_),
    .C(_2876_),
    .Y(_0934_));
 OR3x2_ASAP7_75t_R _6438_ (.A(_0685_),
    .B(_3044_),
    .C(_3046_),
    .Y(_3058_));
 AO32x2_ASAP7_75t_R _6439_ (.A1(_2876_),
    .A2(_3036_),
    .A3(_3058_),
    .B1(_2979_),
    .B2(net31),
    .Y(_0935_));
 AND2x2_ASAP7_75t_R _6440_ (.A(net32),
    .B(_2827_),
    .Y(_3059_));
 XNOR2x2_ASAP7_75t_R _6441_ (.A(_0857_),
    .B(_0684_),
    .Y(_3060_));
 OR2x2_ASAP7_75t_R _6442_ (.A(_3059_),
    .B(_3060_),
    .Y(_3061_));
 OA221x2_ASAP7_75t_R _6443_ (.A1(_3036_),
    .A2(_3059_),
    .B1(_3061_),
    .B2(_3056_),
    .C(_2876_),
    .Y(_0936_));
 OR3x2_ASAP7_75t_R _6444_ (.A(_0687_),
    .B(_3044_),
    .C(_3046_),
    .Y(_3062_));
 AO32x2_ASAP7_75t_R _6445_ (.A1(_2876_),
    .A2(_3036_),
    .A3(_3062_),
    .B1(_2979_),
    .B2(net33),
    .Y(_0937_));
 AND2x2_ASAP7_75t_R _6446_ (.A(net34),
    .B(_2827_),
    .Y(_3063_));
 XNOR2x2_ASAP7_75t_R _6447_ (.A(_0855_),
    .B(_0686_),
    .Y(_3064_));
 OR2x2_ASAP7_75t_R _6448_ (.A(_3063_),
    .B(_3064_),
    .Y(_3065_));
 OA221x2_ASAP7_75t_R _6449_ (.A1(_3036_),
    .A2(_3063_),
    .B1(_3065_),
    .B2(_3056_),
    .C(_2876_),
    .Y(_0938_));
 OR3x2_ASAP7_75t_R _6450_ (.A(_0689_),
    .B(_3044_),
    .C(_3046_),
    .Y(_3066_));
 AO32x2_ASAP7_75t_R _6451_ (.A1(_2876_),
    .A2(_3036_),
    .A3(_3066_),
    .B1(_2979_),
    .B2(net35),
    .Y(_0939_));
 AND2x2_ASAP7_75t_R _6452_ (.A(net36),
    .B(_2827_),
    .Y(_3067_));
 XNOR2x2_ASAP7_75t_R _6453_ (.A(_0853_),
    .B(_0688_),
    .Y(_3068_));
 OR2x2_ASAP7_75t_R _6454_ (.A(_3067_),
    .B(_3068_),
    .Y(_3069_));
 OA221x2_ASAP7_75t_R _6455_ (.A1(_3036_),
    .A2(_3067_),
    .B1(_3069_),
    .B2(_3056_),
    .C(_2876_),
    .Y(_0940_));
 OR3x2_ASAP7_75t_R _6456_ (.A(_0691_),
    .B(_3044_),
    .C(_3046_),
    .Y(_3070_));
 AO32x2_ASAP7_75t_R _6457_ (.A1(_2876_),
    .A2(_3036_),
    .A3(_3070_),
    .B1(_2979_),
    .B2(net22),
    .Y(_0941_));
 AND2x2_ASAP7_75t_R _6458_ (.A(net23),
    .B(_2827_),
    .Y(_3071_));
 XNOR2x2_ASAP7_75t_R _6459_ (.A(_0690_),
    .B(_0851_),
    .Y(_3072_));
 OR2x2_ASAP7_75t_R _6460_ (.A(_3071_),
    .B(_3072_),
    .Y(_3073_));
 OA221x2_ASAP7_75t_R _6461_ (.A1(_3036_),
    .A2(_3071_),
    .B1(_3073_),
    .B2(_3056_),
    .C(_2876_),
    .Y(_0942_));
 OR3x2_ASAP7_75t_R _6462_ (.A(_0693_),
    .B(_3044_),
    .C(_3046_),
    .Y(_3074_));
 AO32x2_ASAP7_75t_R _6463_ (.A1(_2876_),
    .A2(_3036_),
    .A3(_3074_),
    .B1(_2979_),
    .B2(net24),
    .Y(_0943_));
 AND2x2_ASAP7_75t_R _6464_ (.A(net25),
    .B(_2827_),
    .Y(_3075_));
 XNOR2x2_ASAP7_75t_R _6465_ (.A(_0692_),
    .B(_0848_),
    .Y(_3076_));
 OR2x2_ASAP7_75t_R _6466_ (.A(_3075_),
    .B(_3076_),
    .Y(_3077_));
 OA221x2_ASAP7_75t_R _6467_ (.A1(_3036_),
    .A2(_3075_),
    .B1(_3077_),
    .B2(_3056_),
    .C(_2876_),
    .Y(_0944_));
 OR3x2_ASAP7_75t_R _6468_ (.A(_0695_),
    .B(_3044_),
    .C(_3046_),
    .Y(_3078_));
 AO32x2_ASAP7_75t_R _6469_ (.A1(_2876_),
    .A2(_3036_),
    .A3(_3078_),
    .B1(_2979_),
    .B2(net26),
    .Y(_0945_));
 XNOR2x2_ASAP7_75t_R _6470_ (.A(_3357_),
    .B(_3018_),
    .Y(_3079_));
 TAPCELL_ASAP7_75t_R PHY_20 ();
 OR2x2_ASAP7_75t_R _6472_ (.A(net27),
    .B(_2831_),
    .Y(_3081_));
 TAPCELL_ASAP7_75t_R PHY_19 ();
 OA211x2_ASAP7_75t_R _6474_ (.A1(_2827_),
    .A2(_3079_),
    .B(_3081_),
    .C(_2876_),
    .Y(_0946_));
 OR2x2_ASAP7_75t_R _6475_ (.A(\__st_3[16] ),
    .B(_2831_),
    .Y(_3083_));
 OA211x2_ASAP7_75t_R _6476_ (.A1(_2827_),
    .A2(_3079_),
    .B(_3083_),
    .C(_2876_),
    .Y(_0947_));
 OR2x2_ASAP7_75t_R _6477_ (.A(\__st_3[17] ),
    .B(_2831_),
    .Y(_3084_));
 OA211x2_ASAP7_75t_R _6478_ (.A1(_2827_),
    .A2(_3079_),
    .B(_3084_),
    .C(_2876_),
    .Y(_0948_));
 OR2x2_ASAP7_75t_R _6479_ (.A(\__st_3[18] ),
    .B(_2831_),
    .Y(_3085_));
 OA211x2_ASAP7_75t_R _6480_ (.A1(_2827_),
    .A2(_3079_),
    .B(_3085_),
    .C(_2876_),
    .Y(_0949_));
 OR2x2_ASAP7_75t_R _6481_ (.A(\__st_3[19] ),
    .B(_2831_),
    .Y(_3086_));
 OA211x2_ASAP7_75t_R _6482_ (.A1(_2827_),
    .A2(_3079_),
    .B(_3086_),
    .C(_2876_),
    .Y(_0950_));
 OR2x2_ASAP7_75t_R _6483_ (.A(\__st_3[20] ),
    .B(_2831_),
    .Y(_3087_));
 OA211x2_ASAP7_75t_R _6484_ (.A1(_2827_),
    .A2(_3079_),
    .B(_3087_),
    .C(_2876_),
    .Y(_0951_));
 OR2x2_ASAP7_75t_R _6485_ (.A(\__st_3[21] ),
    .B(_2831_),
    .Y(_3088_));
 OA211x2_ASAP7_75t_R _6486_ (.A1(_2827_),
    .A2(_3079_),
    .B(_3088_),
    .C(_2876_),
    .Y(_0952_));
 OR2x2_ASAP7_75t_R _6487_ (.A(\__st_3[22] ),
    .B(_2831_),
    .Y(_3089_));
 OA211x2_ASAP7_75t_R _6488_ (.A1(_2827_),
    .A2(_3079_),
    .B(_3089_),
    .C(_2876_),
    .Y(_0953_));
 OR2x2_ASAP7_75t_R _6489_ (.A(\__st_3[23] ),
    .B(_2831_),
    .Y(_3090_));
 OA211x2_ASAP7_75t_R _6490_ (.A1(_2827_),
    .A2(_3079_),
    .B(_3090_),
    .C(_2876_),
    .Y(_0954_));
 OR2x2_ASAP7_75t_R _6491_ (.A(\__st_3[24] ),
    .B(_2831_),
    .Y(_3091_));
 OA211x2_ASAP7_75t_R _6492_ (.A1(_2827_),
    .A2(_3079_),
    .B(_3091_),
    .C(_2876_),
    .Y(_0955_));
 OR2x2_ASAP7_75t_R _6493_ (.A(\__st_3[25] ),
    .B(_2831_),
    .Y(_3092_));
 TAPCELL_ASAP7_75t_R PHY_18 ();
 OA211x2_ASAP7_75t_R _6495_ (.A1(_2827_),
    .A2(_3079_),
    .B(_3092_),
    .C(_2876_),
    .Y(_0956_));
 OR2x2_ASAP7_75t_R _6496_ (.A(\__st_3[26] ),
    .B(_2831_),
    .Y(_3094_));
 OA211x2_ASAP7_75t_R _6497_ (.A1(_2827_),
    .A2(_3079_),
    .B(_3094_),
    .C(_2876_),
    .Y(_0957_));
 OR2x2_ASAP7_75t_R _6498_ (.A(\__st_3[27] ),
    .B(_2831_),
    .Y(_3095_));
 OA211x2_ASAP7_75t_R _6499_ (.A1(_2827_),
    .A2(_3079_),
    .B(_3095_),
    .C(_2876_),
    .Y(_0958_));
 OR2x2_ASAP7_75t_R _6500_ (.A(\__st_3[28] ),
    .B(_2831_),
    .Y(_3096_));
 OA211x2_ASAP7_75t_R _6501_ (.A1(_2827_),
    .A2(_3079_),
    .B(_3096_),
    .C(_2876_),
    .Y(_0959_));
 OR2x2_ASAP7_75t_R _6502_ (.A(\__st_3[29] ),
    .B(_2831_),
    .Y(_3097_));
 OA211x2_ASAP7_75t_R _6503_ (.A1(_2827_),
    .A2(_3079_),
    .B(_3097_),
    .C(_2876_),
    .Y(_0960_));
 INVx2_ASAP7_75t_R _6504_ (.A(_3356_),
    .Y(_3098_));
 OR2x2_ASAP7_75t_R _6505_ (.A(_3098_),
    .B(_2831_),
    .Y(_3099_));
 OA211x2_ASAP7_75t_R _6506_ (.A1(_2827_),
    .A2(_3079_),
    .B(_3099_),
    .C(_2876_),
    .Y(_0961_));
 INVx2_ASAP7_75t_R _6507_ (.A(_0529_),
    .Y(_3100_));
 OR2x2_ASAP7_75t_R _6508_ (.A(_3100_),
    .B(_2831_),
    .Y(_3101_));
 OA211x2_ASAP7_75t_R _6509_ (.A1(_2827_),
    .A2(_3079_),
    .B(_3101_),
    .C(_2876_),
    .Y(_0962_));
 TAPCELL_ASAP7_75t_R PHY_17 ();
 INVx2_ASAP7_75t_R _6511_ (.A(_3405_),
    .Y(_3103_));
 OR2x2_ASAP7_75t_R _6512_ (.A(_3103_),
    .B(net20),
    .Y(_3104_));
 OA211x2_ASAP7_75t_R _6513_ (.A1(net1),
    .A2(_2756_),
    .B(_3104_),
    .C(_2876_),
    .Y(_0963_));
 OR2x2_ASAP7_75t_R _6514_ (.A(\__in_sample_reg[1] ),
    .B(net20),
    .Y(_3105_));
 OA211x2_ASAP7_75t_R _6515_ (.A1(net8),
    .A2(_2756_),
    .B(_3105_),
    .C(_2876_),
    .Y(_0964_));
 OR2x2_ASAP7_75t_R _6516_ (.A(\__in_sample_reg[2] ),
    .B(net20),
    .Y(_3106_));
 OA211x2_ASAP7_75t_R _6517_ (.A1(net9),
    .A2(_2756_),
    .B(_3106_),
    .C(_2876_),
    .Y(_0965_));
 OR2x2_ASAP7_75t_R _6518_ (.A(\__in_sample_reg[3] ),
    .B(net20),
    .Y(_3107_));
 TAPCELL_ASAP7_75t_R PHY_16 ();
 OA211x2_ASAP7_75t_R _6520_ (.A1(net10),
    .A2(_2756_),
    .B(_3107_),
    .C(_2876_),
    .Y(_0966_));
 OR2x2_ASAP7_75t_R _6521_ (.A(\__in_sample_reg[4] ),
    .B(net20),
    .Y(_3109_));
 OA211x2_ASAP7_75t_R _6522_ (.A1(net11),
    .A2(_2756_),
    .B(_3109_),
    .C(_2876_),
    .Y(_0967_));
 OR2x2_ASAP7_75t_R _6523_ (.A(\__in_sample_reg[5] ),
    .B(net20),
    .Y(_3110_));
 OA211x2_ASAP7_75t_R _6524_ (.A1(net12),
    .A2(_2756_),
    .B(_3110_),
    .C(_2876_),
    .Y(_0968_));
 OR2x2_ASAP7_75t_R _6525_ (.A(\__in_sample_reg[6] ),
    .B(net20),
    .Y(_3111_));
 OA211x2_ASAP7_75t_R _6526_ (.A1(net13),
    .A2(_2756_),
    .B(_3111_),
    .C(_2876_),
    .Y(_0969_));
 OR2x2_ASAP7_75t_R _6527_ (.A(\__in_sample_reg[7] ),
    .B(net20),
    .Y(_3112_));
 OA211x2_ASAP7_75t_R _6528_ (.A1(net14),
    .A2(_2756_),
    .B(_3112_),
    .C(_2876_),
    .Y(_0970_));
 OR2x2_ASAP7_75t_R _6529_ (.A(\__in_sample_reg[8] ),
    .B(net20),
    .Y(_3113_));
 OA211x2_ASAP7_75t_R _6530_ (.A1(net15),
    .A2(_2756_),
    .B(_3113_),
    .C(_2876_),
    .Y(_0971_));
 OR2x2_ASAP7_75t_R _6531_ (.A(\__in_sample_reg[9] ),
    .B(net20),
    .Y(_3114_));
 OA211x2_ASAP7_75t_R _6532_ (.A1(net16),
    .A2(_2756_),
    .B(_3114_),
    .C(_2876_),
    .Y(_0972_));
 OR2x2_ASAP7_75t_R _6533_ (.A(\__in_sample_reg[10] ),
    .B(net20),
    .Y(_3115_));
 OA211x2_ASAP7_75t_R _6534_ (.A1(net2),
    .A2(_2756_),
    .B(_3115_),
    .C(_2876_),
    .Y(_0973_));
 OR2x2_ASAP7_75t_R _6535_ (.A(\__in_sample_reg[11] ),
    .B(net20),
    .Y(_3116_));
 OA211x2_ASAP7_75t_R _6536_ (.A1(net3),
    .A2(_2756_),
    .B(_3116_),
    .C(_2876_),
    .Y(_0974_));
 OR2x2_ASAP7_75t_R _6537_ (.A(\__in_sample_reg[12] ),
    .B(net20),
    .Y(_3117_));
 OA211x2_ASAP7_75t_R _6538_ (.A1(net4),
    .A2(_2756_),
    .B(_3117_),
    .C(_2876_),
    .Y(_0975_));
 OR2x2_ASAP7_75t_R _6539_ (.A(\__in_sample_reg[13] ),
    .B(net20),
    .Y(_3118_));
 OA211x2_ASAP7_75t_R _6540_ (.A1(net5),
    .A2(_2756_),
    .B(_3118_),
    .C(_2876_),
    .Y(_0976_));
 OR2x2_ASAP7_75t_R _6541_ (.A(\__in_sample_reg[14] ),
    .B(net20),
    .Y(_3119_));
 OA211x2_ASAP7_75t_R _6542_ (.A1(net6),
    .A2(_2756_),
    .B(_3119_),
    .C(_2876_),
    .Y(_0977_));
 OR2x2_ASAP7_75t_R _6543_ (.A(\__in_sample_reg[15] ),
    .B(net20),
    .Y(_3120_));
 OA211x2_ASAP7_75t_R _6544_ (.A1(net7),
    .A2(_2756_),
    .B(_3120_),
    .C(_2876_),
    .Y(_0978_));
 INVx2_ASAP7_75t_R _6545_ (.A(_2755_),
    .Y(_3121_));
 OA21x2_ASAP7_75t_R _6546_ (.A1(net17),
    .A2(_3121_),
    .B(_2876_),
    .Y(_0979_));
 AO21x2_ASAP7_75t_R _6547_ (.A1(_0427_),
    .A2(_2754_),
    .B(net19),
    .Y(_3122_));
 INVx2_ASAP7_75t_R _6548_ (.A(_3122_),
    .Y(_0980_));
 INVx2_ASAP7_75t_R _6549_ (.A(_0768_),
    .Y(_3235_));
 INVx2_ASAP7_75t_R _6550_ (.A(_0769_),
    .Y(_3253_));
 INVx2_ASAP7_75t_R _6551_ (.A(_3646_),
    .Y(_3269_));
 INVx2_ASAP7_75t_R _6552_ (.A(_0012_),
    .Y(_3173_));
 INVx2_ASAP7_75t_R _6553_ (.A(_0812_),
    .Y(_3294_));
 INVx2_ASAP7_75t_R _6554_ (.A(_0845_),
    .Y(_3355_));
 INVx2_ASAP7_75t_R _6555_ (.A(_3720_),
    .Y(_3375_));
 INVx2_ASAP7_75t_R _6556_ (.A(_0059_),
    .Y(_3179_));
 INVx2_ASAP7_75t_R _6557_ (.A(net238),
    .Y(_3125_));
 INVx2_ASAP7_75t_R _6558_ (.A(_0729_),
    .Y(_3210_));
 INVx2_ASAP7_75t_R _6559_ (.A(_0767_),
    .Y(_3219_));
 FAx1_ASAP7_75t_R _6560_ (.SN(_0452_),
    .A(_3123_),
    .B(\__in_sample_reg[1] ),
    .CI(_3124_),
    .CON(_0452_));
 FAx1_ASAP7_75t_R _6561_ (.SN(_3433_),
    .A(_3126_),
    .B(\__in_sample_reg[2] ),
    .CI(_3125_),
    .CON(_0455_));
 FAx1_ASAP7_75t_R _6562_ (.SN(_3440_),
    .A(_3127_),
    .B(\__in_sample_reg[6] ),
    .CI(_3128_),
    .CON(_0460_));
 FAx1_ASAP7_75t_R _6563_ (.SN(_3449_),
    .A(\__st_1[4] ),
    .B(_3129_),
    .CI(_3130_),
    .CON(_0461_));
 FAx1_ASAP7_75t_R _6564_ (.SN(_3453_),
    .A(_3131_),
    .B(\__in_sample_reg[14] ),
    .CI(_3132_),
    .CON(_0468_));
 FAx1_ASAP7_75t_R _6565_ (.SN(_3459_),
    .A(_3133_),
    .B(\__in_sample_reg[12] ),
    .CI(_3134_),
    .CON(_0469_));
 FAx1_ASAP7_75t_R _6566_ (.SN(_3466_),
    .A(_3135_),
    .B(\__in_sample_reg[10] ),
    .CI(_3136_),
    .CON(_0470_));
 FAx1_ASAP7_75t_R _6567_ (.SN(_3475_),
    .A(_3137_),
    .B(\__in_sample_reg[8] ),
    .CI(_3138_),
    .CON(_0471_));
 FAx1_ASAP7_75t_R _6568_ (.SN(_3479_),
    .A(_3139_),
    .B(\__in_sample_reg[15] ),
    .CI(_3140_),
    .CON(_0453_));
 FAx1_ASAP7_75t_R _6569_ (.SN(_3481_),
    .A(_3141_),
    .B(\__in_sample_reg[15] ),
    .CI(_3142_),
    .CON(_0483_));
 FAx1_ASAP7_75t_R _6570_ (.SN(_3483_),
    .A(_3143_),
    .B(\__in_sample_reg[15] ),
    .CI(_3144_),
    .CON(_0484_));
 FAx1_ASAP7_75t_R _6571_ (.SN(_3485_),
    .A(\__st_1[24] ),
    .B(_3145_),
    .CI(_3146_),
    .CON(_0568_));
 FAx1_ASAP7_75t_R _6572_ (.SN(_3487_),
    .A(\__st_1[22] ),
    .B(_3145_),
    .CI(_3147_),
    .CON(_0569_));
 FAx1_ASAP7_75t_R _6573_ (.SN(_3489_),
    .A(\__st_1[20] ),
    .B(_3145_),
    .CI(_3148_),
    .CON(_0570_));
 FAx1_ASAP7_75t_R _6574_ (.SN(_3491_),
    .A(\__st_1[18] ),
    .B(_3145_),
    .CI(_3149_),
    .CON(_0571_));
 FAx1_ASAP7_75t_R _6575_ (.SN(_3493_),
    .A(\__st_1[16] ),
    .B(_3145_),
    .CI(_3150_),
    .CON(_0572_));
 FAx1_ASAP7_75t_R _6576_ (.SN(_0022_),
    .A(_3151_),
    .B(_3152_),
    .CI(_3153_),
    .CON(_0021_));
 FAx1_ASAP7_75t_R _6577_ (.SN(_0026_),
    .A(_3156_),
    .B(_3157_),
    .CI(_3158_),
    .CON(_0023_));
 FAx1_ASAP7_75t_R _6578_ (.SN(_0030_),
    .A(_3159_),
    .B(_3160_),
    .CI(_3161_),
    .CON(_0028_));
 FAx1_ASAP7_75t_R _6579_ (.SN(_0035_),
    .A(_3162_),
    .B(_3163_),
    .CI(_3164_),
    .CON(_0033_));
 FAx1_ASAP7_75t_R _6580_ (.SN(_0040_),
    .A(_3165_),
    .B(_3166_),
    .CI(_3167_),
    .CON(_0038_));
 FAx1_ASAP7_75t_R _6581_ (.SN(_0045_),
    .A(_3168_),
    .B(_3169_),
    .CI(_3170_),
    .CON(_0043_));
 FAx1_ASAP7_75t_R _6582_ (.SN(_0050_),
    .A(_3171_),
    .B(_3172_),
    .CI(_3173_),
    .CON(_0048_));
 FAx1_ASAP7_75t_R _6583_ (.SN(_0053_),
    .A(_3174_),
    .B(_3175_),
    .CI(_3176_),
    .CON(_0012_));
 FAx1_ASAP7_75t_R _6584_ (.SN(_0056_),
    .A(_3171_),
    .B(_3177_),
    .CI(_3178_),
    .CON(_0059_));
 FAx1_ASAP7_75t_R _6585_ (.SN(_0061_),
    .A(_3180_),
    .B(_3181_),
    .CI(_3179_),
    .CON(_0060_));
 FAx1_ASAP7_75t_R _6586_ (.SN(_0068_),
    .A(_3182_),
    .B(_3183_),
    .CI(_3184_),
    .CON(_0067_));
 FAx1_ASAP7_75t_R _6587_ (.SN(_0071_),
    .A(_3185_),
    .B(_3186_),
    .CI(_3187_),
    .CON(_0070_));
 FAx1_ASAP7_75t_R _6588_ (.SN(_0082_),
    .A(_3188_),
    .B(_3189_),
    .CI(_3190_),
    .CON(_0081_));
 FAx1_ASAP7_75t_R _6589_ (.SN(_0574_),
    .A(_3191_),
    .B(_1570_),
    .CI(_3193_),
    .CON(_0573_));
 FAx1_ASAP7_75t_R _6590_ (.SN(_0086_),
    .A(_3194_),
    .B(_3195_),
    .CI(_3196_),
    .CON(_0085_));
 FAx1_ASAP7_75t_R _6591_ (.SN(_0576_),
    .A(_3197_),
    .B(net38),
    .CI(_3199_),
    .CON(_0575_));
 FAx1_ASAP7_75t_R _6592_ (.SN(_0578_),
    .A(_3200_),
    .B(net38),
    .CI(_3201_),
    .CON(_0577_));
 FAx1_ASAP7_75t_R _6593_ (.SN(_0580_),
    .A(_3202_),
    .B(net38),
    .CI(_3203_),
    .CON(_0579_));
 FAx1_ASAP7_75t_R _6594_ (.SN(_0582_),
    .A(\__st_0[8] ),
    .B(net229),
    .CI(_3205_),
    .CON(_0581_));
 FAx1_ASAP7_75t_R _6595_ (.SN(_0584_),
    .A(_3206_),
    .B(_1727_),
    .CI(_3208_),
    .CON(_0583_));
 FAx1_ASAP7_75t_R _6596_ (.SN(_0116_),
    .A(\__st_0[1] ),
    .B(_3209_),
    .CI(_3210_),
    .CON(_3208_));
 FAx1_ASAP7_75t_R _6597_ (.SN(_0586_),
    .A(_3188_),
    .B(_3159_),
    .CI(_3211_),
    .CON(_0585_));
 FAx1_ASAP7_75t_R _6598_ (.SN(_0588_),
    .A(_1363_),
    .B(_3162_),
    .CI(_3213_),
    .CON(_0587_));
 FAx1_ASAP7_75t_R _6599_ (.SN(_0590_),
    .A(_3165_),
    .B(_3194_),
    .CI(_3214_),
    .CON(_0589_));
 FAx1_ASAP7_75t_R _6600_ (.SN(_0592_),
    .A(_3182_),
    .B(_3168_),
    .CI(_3215_),
    .CON(_0591_));
 FAx1_ASAP7_75t_R _6601_ (.SN(_0594_),
    .A(_3171_),
    .B(_3185_),
    .CI(_3216_),
    .CON(_0593_));
 FAx1_ASAP7_75t_R _6602_ (.SN(_0157_),
    .A(_3217_),
    .B(_1336_),
    .CI(_3219_),
    .CON(_3216_));
 FAx1_ASAP7_75t_R _6603_ (.SN(_0160_),
    .A(_1348_),
    .B(_3221_),
    .CI(_3222_),
    .CON(_0159_));
 FAx1_ASAP7_75t_R _6604_ (.SN(_0596_),
    .A(_1363_),
    .B(_3223_),
    .CI(_3224_),
    .CON(_0595_));
 FAx1_ASAP7_75t_R _6605_ (.SN(_0598_),
    .A(_3194_),
    .B(_3225_),
    .CI(_3226_),
    .CON(_0597_));
 FAx1_ASAP7_75t_R _6606_ (.SN(_0600_),
    .A(_3182_),
    .B(_3227_),
    .CI(_3228_),
    .CON(_0599_));
 FAx1_ASAP7_75t_R _6607_ (.SN(_0602_),
    .A(_3185_),
    .B(_3229_),
    .CI(_3230_),
    .CON(_0601_));
 FAx1_ASAP7_75t_R _6608_ (.SN(_0604_),
    .A(_3180_),
    .B(_3231_),
    .CI(_3232_),
    .CON(_0603_));
 FAx1_ASAP7_75t_R _6609_ (.SN(_0178_),
    .A(_3233_),
    .B(_3234_),
    .CI(_3235_),
    .CON(_3232_));
 FAx1_ASAP7_75t_R _6610_ (.SN(_0606_),
    .A(_3151_),
    .B(_3236_),
    .CI(_3237_),
    .CON(_0605_));
 FAx1_ASAP7_75t_R _6611_ (.SN(_0182_),
    .A(_3239_),
    .B(_3240_),
    .CI(_3241_),
    .CON(_0181_));
 FAx1_ASAP7_75t_R _6612_ (.SN(_0183_),
    .A(_3159_),
    .B(_1935_),
    .CI(_3243_),
    .CON(_0607_));
 FAx1_ASAP7_75t_R _6613_ (.SN(_0185_),
    .A(_3244_),
    .B(_3245_),
    .CI(_3246_),
    .CON(_0184_));
 FAx1_ASAP7_75t_R _6614_ (.SN(_0186_),
    .A(_3165_),
    .B(_3247_),
    .CI(_3248_),
    .CON(_0608_));
 FAx1_ASAP7_75t_R _6615_ (.SN(_0187_),
    .A(_3168_),
    .B(_3249_),
    .CI(_3250_),
    .CON(_0609_));
 FAx1_ASAP7_75t_R _6616_ (.SN(_0188_),
    .A(_1207_),
    .B(_3252_),
    .CI(_3253_),
    .CON(_3250_));
 FAx1_ASAP7_75t_R _6617_ (.SN(_0611_),
    .A(_3139_),
    .B(_3254_),
    .CI(_3255_),
    .CON(_0610_));
 FAx1_ASAP7_75t_R _6618_ (.SN(_0613_),
    .A(_3141_),
    .B(_3254_),
    .CI(_3256_),
    .CON(_0612_));
 FAx1_ASAP7_75t_R _6619_ (.SN(_0615_),
    .A(_3143_),
    .B(_3254_),
    .CI(_3257_),
    .CON(_0614_));
 FAx1_ASAP7_75t_R _6620_ (.SN(_0617_),
    .A(_3258_),
    .B(_3254_),
    .CI(_3259_),
    .CON(_0616_));
 FAx1_ASAP7_75t_R _6621_ (.SN(_0619_),
    .A(\__st_1[22] ),
    .B(_3260_),
    .CI(_3261_),
    .CON(_0618_));
 FAx1_ASAP7_75t_R _6622_ (.SN(_0621_),
    .A(_3262_),
    .B(_3254_),
    .CI(_3263_),
    .CON(_0620_));
 FAx1_ASAP7_75t_R _6623_ (.SN(_0623_),
    .A(\__st_1[18] ),
    .B(_3260_),
    .CI(_3264_),
    .CON(_0622_));
 FAx1_ASAP7_75t_R _6624_ (.SN(_0242_),
    .A(_3265_),
    .B(_3266_),
    .CI(_3267_),
    .CON(_0241_));
 FAx1_ASAP7_75t_R _6625_ (.SN(_0624_),
    .A(_3123_),
    .B(_3268_),
    .CI(_3269_),
    .CON(_3647_));
 FAx1_ASAP7_75t_R _6626_ (.SN(_0626_),
    .A(_3126_),
    .B(_3271_),
    .CI(_3270_),
    .CON(_0625_));
 FAx1_ASAP7_75t_R _6627_ (.SN(_0628_),
    .A(_3272_),
    .B(_3273_),
    .CI(_3274_),
    .CON(_0627_));
 FAx1_ASAP7_75t_R _6628_ (.SN(_0630_),
    .A(_3127_),
    .B(_3275_),
    .CI(_3276_),
    .CON(_0629_));
 FAx1_ASAP7_75t_R _6629_ (.SN(_0632_),
    .A(_3137_),
    .B(_3277_),
    .CI(_2137_),
    .CON(_0631_));
 FAx1_ASAP7_75t_R _6630_ (.SN(_0634_),
    .A(_3135_),
    .B(_3279_),
    .CI(_3280_),
    .CON(_0633_));
 FAx1_ASAP7_75t_R _6631_ (.SN(_0636_),
    .A(_3133_),
    .B(_3281_),
    .CI(_3282_),
    .CON(_0635_));
 FAx1_ASAP7_75t_R _6632_ (.SN(_0638_),
    .A(\__st_1[14] ),
    .B(_3283_),
    .CI(_3284_),
    .CON(_0637_));
 FAx1_ASAP7_75t_R _6633_ (.SN(_0640_),
    .A(_3285_),
    .B(net38),
    .CI(_3286_),
    .CON(_0639_));
 FAx1_ASAP7_75t_R _6634_ (.SN(_0642_),
    .A(_3287_),
    .B(net38),
    .CI(_3288_),
    .CON(_0641_));
 FAx1_ASAP7_75t_R _6635_ (.SN(_0644_),
    .A(_3289_),
    .B(net38),
    .CI(_3290_),
    .CON(_0643_));
 FAx1_ASAP7_75t_R _6636_ (.SN(_0646_),
    .A(\__st_2[8] ),
    .B(net229),
    .CI(_3291_),
    .CON(_0645_));
 FAx1_ASAP7_75t_R _6637_ (.SN(_0648_),
    .A(_3292_),
    .B(_1727_),
    .CI(_3293_),
    .CON(_0647_));
 FAx1_ASAP7_75t_R _6638_ (.SN(_0264_),
    .A(\__st_2[1] ),
    .B(_3209_),
    .CI(_3294_),
    .CON(_3293_));
 FAx1_ASAP7_75t_R _6639_ (.SN(_0650_),
    .A(_3295_),
    .B(_3296_),
    .CI(_3297_),
    .CON(_0649_));
 FAx1_ASAP7_75t_R _6640_ (.SN(_0652_),
    .A(_3298_),
    .B(_3299_),
    .CI(_3300_),
    .CON(_0651_));
 FAx1_ASAP7_75t_R _6641_ (.SN(_0654_),
    .A(_3301_),
    .B(_3302_),
    .CI(_3303_),
    .CON(_0653_));
 FAx1_ASAP7_75t_R _6642_ (.SN(_0300_),
    .A(_2333_),
    .B(_2417_),
    .CI(_3306_),
    .CON(_0298_));
 FAx1_ASAP7_75t_R _6643_ (.SN(_0656_),
    .A(_2383_),
    .B(_3308_),
    .CI(_3309_),
    .CON(_0655_));
 FAx1_ASAP7_75t_R _6644_ (.SN(_0657_),
    .A(_3310_),
    .B(_2484_),
    .CI(_3312_),
    .CON(_3667_));
 FAx1_ASAP7_75t_R _6645_ (.SN(_0659_),
    .A(_3295_),
    .B(_2512_),
    .CI(_3314_),
    .CON(_0658_));
 FAx1_ASAP7_75t_R _6646_ (.SN(_0311_),
    .A(_2261_),
    .B(_3318_),
    .CI(_3319_),
    .CON(_0310_));
 FAx1_ASAP7_75t_R _6647_ (.SN(_0316_),
    .A(_2290_),
    .B(_2551_),
    .CI(_3322_),
    .CON(_0314_));
 FAx1_ASAP7_75t_R _6648_ (.SN(_0321_),
    .A(_2333_),
    .B(_2558_),
    .CI(_3324_),
    .CON(_0319_));
 FAx1_ASAP7_75t_R _6649_ (.SN(_0326_),
    .A(_3325_),
    .B(_3326_),
    .CI(_3327_),
    .CON(_0324_));
 FAx1_ASAP7_75t_R _6650_ (.SN(_0661_),
    .A(_3328_),
    .B(_3329_),
    .CI(_3330_),
    .CON(_0660_));
 FAx1_ASAP7_75t_R _6651_ (.SN(_0662_),
    .A(_3308_),
    .B(_3331_),
    .CI(_3332_),
    .CON(_3677_));
 FAx1_ASAP7_75t_R _6652_ (.SN(_0664_),
    .A(_2202_),
    .B(_2529_),
    .CI(_3336_),
    .CON(_0663_));
 FAx1_ASAP7_75t_R _6653_ (.SN(_0334_),
    .A(_2240_),
    .B(_2547_),
    .CI(_3341_),
    .CON(_0333_));
 FAx1_ASAP7_75t_R _6654_ (.SN(_0336_),
    .A(_2271_),
    .B(_2553_),
    .CI(_3344_),
    .CON(_0335_));
 FAx1_ASAP7_75t_R _6655_ (.SN(_0338_),
    .A(_2315_),
    .B(_3346_),
    .CI(_3347_),
    .CON(_0337_));
 FAx1_ASAP7_75t_R _6656_ (.SN(_0340_),
    .A(_3348_),
    .B(_2566_),
    .CI(_3350_),
    .CON(_0339_));
 FAx1_ASAP7_75t_R _6657_ (.SN(_0666_),
    .A(_3310_),
    .B(_2532_),
    .CI(_3352_),
    .CON(_0665_));
 FAx1_ASAP7_75t_R _6658_ (.SN(_0341_),
    .A(_2436_),
    .B(_3354_),
    .CI(_3355_),
    .CON(_3352_));
 FAx1_ASAP7_75t_R _6659_ (.SN(_0668_),
    .A(_3356_),
    .B(_3357_),
    .CI(_3358_),
    .CON(_0667_));
 FAx1_ASAP7_75t_R _6660_ (.SN(_0670_),
    .A(_3359_),
    .B(_3357_),
    .CI(_3360_),
    .CON(_0669_));
 FAx1_ASAP7_75t_R _6661_ (.SN(_0672_),
    .A(_3361_),
    .B(_3357_),
    .CI(_3362_),
    .CON(_0671_));
 FAx1_ASAP7_75t_R _6662_ (.SN(_0674_),
    .A(_3363_),
    .B(_3357_),
    .CI(_3364_),
    .CON(_0673_));
 FAx1_ASAP7_75t_R _6663_ (.SN(_0676_),
    .A(\__st_3[22] ),
    .B(_3365_),
    .CI(_3366_),
    .CON(_0675_));
 FAx1_ASAP7_75t_R _6664_ (.SN(_0678_),
    .A(_3367_),
    .B(_3357_),
    .CI(_3368_),
    .CON(_0677_));
 FAx1_ASAP7_75t_R _6665_ (.SN(_0680_),
    .A(_3369_),
    .B(_3357_),
    .CI(_3370_),
    .CON(_0679_));
 FAx1_ASAP7_75t_R _6666_ (.SN(_0412_),
    .A(\__st_3[16] ),
    .B(_3371_),
    .CI(_3372_),
    .CON(_0411_));
 FAx1_ASAP7_75t_R _6667_ (.SN(_0681_),
    .A(_3373_),
    .B(_3374_),
    .CI(_3375_),
    .CON(_3721_));
 FAx1_ASAP7_75t_R _6668_ (.SN(_0683_),
    .A(_3377_),
    .B(_3378_),
    .CI(_3376_),
    .CON(_0682_));
 FAx1_ASAP7_75t_R _6669_ (.SN(_0685_),
    .A(_3379_),
    .B(_3380_),
    .CI(_3381_),
    .CON(_0684_));
 FAx1_ASAP7_75t_R _6670_ (.SN(_0687_),
    .A(_3382_),
    .B(_3383_),
    .CI(_3384_),
    .CON(_0686_));
 FAx1_ASAP7_75t_R _6671_ (.SN(_0689_),
    .A(_3385_),
    .B(_3386_),
    .CI(_3387_),
    .CON(_0688_));
 FAx1_ASAP7_75t_R _6672_ (.SN(_0691_),
    .A(_3388_),
    .B(_3389_),
    .CI(_3390_),
    .CON(_0690_));
 FAx1_ASAP7_75t_R _6673_ (.SN(_0693_),
    .A(_3391_),
    .B(_3392_),
    .CI(_3393_),
    .CON(_0692_));
 FAx1_ASAP7_75t_R _6674_ (.SN(_0695_),
    .A(_3394_),
    .B(_3395_),
    .CI(_3396_),
    .CON(_0694_));
 HAxp5_ASAP7_75t_R _6675_ (.A(_1034_),
    .B(_3398_),
    .CON(_0243_),
    .SN(_0696_));
 HAxp5_ASAP7_75t_R _6676_ (.A(_3400_),
    .B(_3399_),
    .CON(_0697_),
    .SN(_0263_));
 HAxp5_ASAP7_75t_R _6677_ (.A(_3401_),
    .B(_3402_),
    .CON(_0698_),
    .SN(_0699_));
 HAxp5_ASAP7_75t_R _6678_ (.A(_3403_),
    .B(_3404_),
    .CON(_0700_),
    .SN(_0459_));
 HAxp5_ASAP7_75t_R _6679_ (.A(\__st_1[0] ),
    .B(_3405_),
    .CON(_3124_),
    .SN(_3408_));
 HAxp5_ASAP7_75t_R _6680_ (.A(_3407_),
    .B(_3408_),
    .CON(_0701_),
    .SN(_0285_));
 HAxp5_ASAP7_75t_R _6681_ (.A(_3409_),
    .B(_3406_),
    .CON(_3176_),
    .SN(_3410_));
 HAxp5_ASAP7_75t_R _6682_ (.A(_3411_),
    .B(\__in_sample_reg[15] ),
    .CON(_0350_),
    .SN(_0352_));
 HAxp5_ASAP7_75t_R _6683_ (.A(_3141_),
    .B(\__in_sample_reg[15] ),
    .CON(_0356_),
    .SN(_0366_));
 HAxp5_ASAP7_75t_R _6684_ (.A(_3412_),
    .B(\__in_sample_reg[15] ),
    .CON(_0373_),
    .SN(_0376_));
 HAxp5_ASAP7_75t_R _6685_ (.A(_3143_),
    .B(\__in_sample_reg[15] ),
    .CON(_0377_),
    .SN(_0380_));
 HAxp5_ASAP7_75t_R _6686_ (.A(_3413_),
    .B(\__in_sample_reg[15] ),
    .CON(_0389_),
    .SN(_0392_));
 HAxp5_ASAP7_75t_R _6687_ (.A(_3258_),
    .B(\__in_sample_reg[15] ),
    .CON(_0397_),
    .SN(_0408_));
 HAxp5_ASAP7_75t_R _6688_ (.A(_3414_),
    .B(\__in_sample_reg[15] ),
    .CON(_0409_),
    .SN(_0410_));
 HAxp5_ASAP7_75t_R _6689_ (.A(_3415_),
    .B(\__in_sample_reg[15] ),
    .CON(_0413_),
    .SN(_0415_));
 HAxp5_ASAP7_75t_R _6690_ (.A(_3416_),
    .B(\__in_sample_reg[15] ),
    .CON(_0416_),
    .SN(_0417_));
 HAxp5_ASAP7_75t_R _6691_ (.A(_3262_),
    .B(\__in_sample_reg[15] ),
    .CON(_0418_),
    .SN(_0419_));
 HAxp5_ASAP7_75t_R _6692_ (.A(_3417_),
    .B(\__in_sample_reg[15] ),
    .CON(_0420_),
    .SN(_0421_));
 HAxp5_ASAP7_75t_R _6693_ (.A(_3418_),
    .B(\__in_sample_reg[15] ),
    .CON(_0422_),
    .SN(_0423_));
 HAxp5_ASAP7_75t_R _6694_ (.A(_3419_),
    .B(\__in_sample_reg[15] ),
    .CON(_0424_),
    .SN(_0425_));
 HAxp5_ASAP7_75t_R _6695_ (.A(_3265_),
    .B(\__in_sample_reg[15] ),
    .CON(_0426_),
    .SN(_0428_));
 HAxp5_ASAP7_75t_R _6696_ (.A(_3420_),
    .B(\__in_sample_reg[15] ),
    .CON(_0429_),
    .SN(_0430_));
 HAxp5_ASAP7_75t_R _6697_ (.A(_3131_),
    .B(\__in_sample_reg[14] ),
    .CON(_0431_),
    .SN(_0432_));
 HAxp5_ASAP7_75t_R _6698_ (.A(_3421_),
    .B(\__in_sample_reg[13] ),
    .CON(_0433_),
    .SN(_0702_));
 HAxp5_ASAP7_75t_R _6699_ (.A(_3133_),
    .B(\__in_sample_reg[12] ),
    .CON(_0434_),
    .SN(_0435_));
 HAxp5_ASAP7_75t_R _6700_ (.A(_3422_),
    .B(\__in_sample_reg[11] ),
    .CON(_0436_),
    .SN(_0703_));
 HAxp5_ASAP7_75t_R _6701_ (.A(_3135_),
    .B(\__in_sample_reg[10] ),
    .CON(_0437_),
    .SN(_0438_));
 HAxp5_ASAP7_75t_R _6702_ (.A(_3423_),
    .B(\__in_sample_reg[9] ),
    .CON(_0439_),
    .SN(_0704_));
 HAxp5_ASAP7_75t_R _6703_ (.A(_3137_),
    .B(\__in_sample_reg[8] ),
    .CON(_0440_),
    .SN(_0441_));
 HAxp5_ASAP7_75t_R _6704_ (.A(_3424_),
    .B(\__in_sample_reg[7] ),
    .CON(_0442_),
    .SN(_0705_));
 HAxp5_ASAP7_75t_R _6705_ (.A(_3127_),
    .B(\__in_sample_reg[6] ),
    .CON(_0443_),
    .SN(_0444_));
 HAxp5_ASAP7_75t_R _6706_ (.A(_3425_),
    .B(\__in_sample_reg[5] ),
    .CON(_0445_),
    .SN(_0446_));
 HAxp5_ASAP7_75t_R _6707_ (.A(_3272_),
    .B(\__in_sample_reg[4] ),
    .CON(_0447_),
    .SN(_0448_));
 HAxp5_ASAP7_75t_R _6708_ (.A(_3426_),
    .B(\__in_sample_reg[3] ),
    .CON(_0449_),
    .SN(_0706_));
 HAxp5_ASAP7_75t_R _6709_ (.A(_3126_),
    .B(\__in_sample_reg[2] ),
    .CON(_0450_),
    .SN(_0451_));
 HAxp5_ASAP7_75t_R _6710_ (.A(_3406_),
    .B(_3427_),
    .CON(_0707_),
    .SN(_0454_));
 HAxp5_ASAP7_75t_R _6711_ (.A(_3217_),
    .B(_1183_),
    .CON(_0502_),
    .SN(_0708_));
 HAxp5_ASAP7_75t_R _6712_ (.A(_1207_),
    .B(_3430_),
    .CON(_0500_),
    .SN(_0709_));
 HAxp5_ASAP7_75t_R _6713_ (.A(_3180_),
    .B(_3431_),
    .CON(_0010_),
    .SN(_3432_));
 HAxp5_ASAP7_75t_R _6714_ (.A(_3433_),
    .B(_3428_),
    .CON(_0456_),
    .SN(_0457_));
 HAxp5_ASAP7_75t_R _6715_ (.A(_3233_),
    .B(_1238_),
    .CON(_0501_),
    .SN(_0458_));
 HAxp5_ASAP7_75t_R _6716_ (.A(_3171_),
    .B(_3172_),
    .CON(_0011_),
    .SN(_3435_));
 HAxp5_ASAP7_75t_R _6717_ (.A(_3436_),
    .B(_3437_),
    .CON(_0496_),
    .SN(_0710_));
 HAxp5_ASAP7_75t_R _6718_ (.A(_3182_),
    .B(_3438_),
    .CON(_0006_),
    .SN(_3439_));
 HAxp5_ASAP7_75t_R _6719_ (.A(_3440_),
    .B(_3441_),
    .CON(_0462_),
    .SN(_0463_));
 HAxp5_ASAP7_75t_R _6720_ (.A(_3442_),
    .B(_1293_),
    .CON(_0497_),
    .SN(_0464_));
 HAxp5_ASAP7_75t_R _6721_ (.A(_3165_),
    .B(_3166_),
    .CON(_0007_),
    .SN(_3444_));
 HAxp5_ASAP7_75t_R _6722_ (.A(_1314_),
    .B(_3446_),
    .CON(_0498_),
    .SN(_0711_));
 HAxp5_ASAP7_75t_R _6723_ (.A(_3185_),
    .B(_3447_),
    .CON(_0008_),
    .SN(_3448_));
 HAxp5_ASAP7_75t_R _6724_ (.A(_3449_),
    .B(_3450_),
    .CON(_0465_),
    .SN(_0466_));
 HAxp5_ASAP7_75t_R _6725_ (.A(_1336_),
    .B(_1338_),
    .CON(_0499_),
    .SN(_0467_));
 HAxp5_ASAP7_75t_R _6726_ (.A(_3168_),
    .B(_3169_),
    .CON(_0009_),
    .SN(_3452_));
 HAxp5_ASAP7_75t_R _6727_ (.A(_3453_),
    .B(_3454_),
    .CON(_0712_),
    .SN(_0472_));
 HAxp5_ASAP7_75t_R _6728_ (.A(_3151_),
    .B(_3152_),
    .CON(_0713_),
    .SN(_0473_));
 HAxp5_ASAP7_75t_R _6729_ (.A(_3154_),
    .B(_3155_),
    .CON(_0489_),
    .SN(_3455_));
 HAxp5_ASAP7_75t_R _6730_ (.A(_1348_),
    .B(_3456_),
    .CON(_0490_),
    .SN(_0714_));
 HAxp5_ASAP7_75t_R _6731_ (.A(_3188_),
    .B(_3457_),
    .CON(_0000_),
    .SN(_3458_));
 HAxp5_ASAP7_75t_R _6732_ (.A(_3459_),
    .B(_3460_),
    .CON(_0474_),
    .SN(_0475_));
 HAxp5_ASAP7_75t_R _6733_ (.A(_3239_),
    .B(_1355_),
    .CON(_0491_),
    .SN(_0476_));
 HAxp5_ASAP7_75t_R _6734_ (.A(_3156_),
    .B(_3157_),
    .CON(_0001_),
    .SN(_3462_));
 HAxp5_ASAP7_75t_R _6735_ (.A(_3191_),
    .B(_3463_),
    .CON(_0492_),
    .SN(_0715_));
 HAxp5_ASAP7_75t_R _6736_ (.A(_1363_),
    .B(_3464_),
    .CON(_0002_),
    .SN(_3465_));
 HAxp5_ASAP7_75t_R _6737_ (.A(_3466_),
    .B(_3467_),
    .CON(_0477_),
    .SN(_0478_));
 HAxp5_ASAP7_75t_R _6738_ (.A(_3468_),
    .B(_1375_),
    .CON(_0493_),
    .SN(_0479_));
 HAxp5_ASAP7_75t_R _6739_ (.A(_3159_),
    .B(_3160_),
    .CON(_0003_),
    .SN(_3470_));
 HAxp5_ASAP7_75t_R _6740_ (.A(_1388_),
    .B(_3472_),
    .CON(_0494_),
    .SN(_0716_));
 HAxp5_ASAP7_75t_R _6741_ (.A(_3194_),
    .B(_3473_),
    .CON(_0004_),
    .SN(_3474_));
 HAxp5_ASAP7_75t_R _6742_ (.A(_3475_),
    .B(_3476_),
    .CON(_0480_),
    .SN(_0481_));
 HAxp5_ASAP7_75t_R _6743_ (.A(_3244_),
    .B(_1402_),
    .CON(_0495_),
    .SN(_0482_));
 HAxp5_ASAP7_75t_R _6744_ (.A(_3162_),
    .B(_3163_),
    .CON(_0005_),
    .SN(_3478_));
 HAxp5_ASAP7_75t_R _6745_ (.A(_3479_),
    .B(_3480_),
    .CON(_0485_),
    .SN(_0717_));
 HAxp5_ASAP7_75t_R _6746_ (.A(_3481_),
    .B(_3482_),
    .CON(_0718_),
    .SN(_0719_));
 HAxp5_ASAP7_75t_R _6747_ (.A(_3483_),
    .B(_3484_),
    .CON(_0486_),
    .SN(_0720_));
 HAxp5_ASAP7_75t_R _6748_ (.A(_3485_),
    .B(_3486_),
    .CON(_0721_),
    .SN(_0722_));
 HAxp5_ASAP7_75t_R _6749_ (.A(_3487_),
    .B(_3488_),
    .CON(_0723_),
    .SN(_0724_));
 HAxp5_ASAP7_75t_R _6750_ (.A(_3489_),
    .B(_3490_),
    .CON(_0487_),
    .SN(_0725_));
 HAxp5_ASAP7_75t_R _6751_ (.A(_3491_),
    .B(_3492_),
    .CON(_0726_),
    .SN(_0727_));
 HAxp5_ASAP7_75t_R _6752_ (.A(_3493_),
    .B(_3494_),
    .CON(_0488_),
    .SN(_0728_));
 HAxp5_ASAP7_75t_R _6753_ (.A(\__st_0[0] ),
    .B(net229),
    .CON(_0729_),
    .SN(_0730_));
 HAxp5_ASAP7_75t_R _6754_ (.A(\__st_0[13] ),
    .B(net229),
    .CON(_0503_),
    .SN(_0731_));
 HAxp5_ASAP7_75t_R _6755_ (.A(\__st_0[12] ),
    .B(net229),
    .CON(_0504_),
    .SN(_0505_));
 HAxp5_ASAP7_75t_R _6756_ (.A(\__st_0[11] ),
    .B(net229),
    .CON(_0506_),
    .SN(_0732_));
 HAxp5_ASAP7_75t_R _6757_ (.A(\__st_0[10] ),
    .B(net229),
    .CON(_0507_),
    .SN(_0508_));
 HAxp5_ASAP7_75t_R _6758_ (.A(\__st_0[9] ),
    .B(net229),
    .CON(_0509_),
    .SN(_0510_));
 HAxp5_ASAP7_75t_R _6759_ (.A(\__st_0[8] ),
    .B(net229),
    .CON(_0511_),
    .SN(_0512_));
 HAxp5_ASAP7_75t_R _6760_ (.A(\__st_0[7] ),
    .B(net229),
    .CON(_0513_),
    .SN(_0514_));
 HAxp5_ASAP7_75t_R _6761_ (.A(_3495_),
    .B(_3496_),
    .CON(_0733_),
    .SN(_0013_));
 HAxp5_ASAP7_75t_R _6762_ (.A(_3497_),
    .B(_3498_),
    .CON(_0734_),
    .SN(_0014_));
 HAxp5_ASAP7_75t_R _6763_ (.A(_3499_),
    .B(_3500_),
    .CON(_0735_),
    .SN(_0015_));
 HAxp5_ASAP7_75t_R _6764_ (.A(_3501_),
    .B(_3502_),
    .CON(_0736_),
    .SN(_0016_));
 HAxp5_ASAP7_75t_R _6765_ (.A(_1532_),
    .B(_3504_),
    .CON(_0737_),
    .SN(_0017_));
 HAxp5_ASAP7_75t_R _6766_ (.A(_3505_),
    .B(_3506_),
    .CON(_0738_),
    .SN(_0018_));
 HAxp5_ASAP7_75t_R _6767_ (.A(_3507_),
    .B(_3508_),
    .CON(_0739_),
    .SN(_0019_));
 HAxp5_ASAP7_75t_R _6768_ (.A(_3509_),
    .B(_3510_),
    .CON(_0740_),
    .SN(_0020_));
 HAxp5_ASAP7_75t_R _6769_ (.A(_3151_),
    .B(_3511_),
    .CON(_0073_),
    .SN(_0025_));
 HAxp5_ASAP7_75t_R _6770_ (.A(_3154_),
    .B(_3512_),
    .CON(_0024_),
    .SN(_3513_));
 HAxp5_ASAP7_75t_R _6771_ (.A(_1348_),
    .B(_1564_),
    .CON(_0741_),
    .SN(_0027_));
 HAxp5_ASAP7_75t_R _6772_ (.A(_3188_),
    .B(_3189_),
    .CON(_0074_),
    .SN(_3515_));
 HAxp5_ASAP7_75t_R _6773_ (.A(_3239_),
    .B(_1568_),
    .CON(_0029_),
    .SN(_0742_));
 HAxp5_ASAP7_75t_R _6774_ (.A(_3156_),
    .B(_3517_),
    .CON(_0075_),
    .SN(_3518_));
 HAxp5_ASAP7_75t_R _6775_ (.A(_3191_),
    .B(_1570_),
    .CON(_0031_),
    .SN(_0032_));
 HAxp5_ASAP7_75t_R _6776_ (.A(_1363_),
    .B(_3519_),
    .CON(_0076_),
    .SN(_3520_));
 HAxp5_ASAP7_75t_R _6777_ (.A(_3468_),
    .B(_1573_),
    .CON(_0034_),
    .SN(_0743_));
 HAxp5_ASAP7_75t_R _6778_ (.A(_3159_),
    .B(_3522_),
    .CON(_0077_),
    .SN(_3523_));
 HAxp5_ASAP7_75t_R _6779_ (.A(_1388_),
    .B(_1575_),
    .CON(_0036_),
    .SN(_0037_));
 HAxp5_ASAP7_75t_R _6780_ (.A(_3194_),
    .B(_3195_),
    .CON(_0078_),
    .SN(_3525_));
 HAxp5_ASAP7_75t_R _6781_ (.A(_3244_),
    .B(_1578_),
    .CON(_0039_),
    .SN(_0744_));
 HAxp5_ASAP7_75t_R _6782_ (.A(_3162_),
    .B(_3527_),
    .CON(_0079_),
    .SN(_3528_));
 HAxp5_ASAP7_75t_R _6783_ (.A(_3436_),
    .B(_1580_),
    .CON(_0041_),
    .SN(_0042_));
 HAxp5_ASAP7_75t_R _6784_ (.A(_3182_),
    .B(_3183_),
    .CON(_0063_),
    .SN(_3530_));
 HAxp5_ASAP7_75t_R _6785_ (.A(_3442_),
    .B(_1583_),
    .CON(_0044_),
    .SN(_0745_));
 HAxp5_ASAP7_75t_R _6786_ (.A(_3165_),
    .B(_3532_),
    .CON(_0064_),
    .SN(_3533_));
 HAxp5_ASAP7_75t_R _6787_ (.A(_1314_),
    .B(_1585_),
    .CON(_0046_),
    .SN(_0047_));
 HAxp5_ASAP7_75t_R _6788_ (.A(_3185_),
    .B(_3186_),
    .CON(_0065_),
    .SN(_3535_));
 HAxp5_ASAP7_75t_R _6789_ (.A(_1336_),
    .B(_1588_),
    .CON(_0049_),
    .SN(_0746_));
 HAxp5_ASAP7_75t_R _6790_ (.A(_3168_),
    .B(_3537_),
    .CON(_0066_),
    .SN(_3538_));
 HAxp5_ASAP7_75t_R _6791_ (.A(_1207_),
    .B(_1590_),
    .CON(_0051_),
    .SN(_0052_));
 HAxp5_ASAP7_75t_R _6792_ (.A(_3180_),
    .B(_3181_),
    .CON(_0058_),
    .SN(_3540_));
 HAxp5_ASAP7_75t_R _6793_ (.A(_3233_),
    .B(_1592_),
    .CON(_0054_),
    .SN(_0747_));
 HAxp5_ASAP7_75t_R _6794_ (.A(_3217_),
    .B(_3542_),
    .CON(_3178_),
    .SN(_0748_));
 HAxp5_ASAP7_75t_R _6795_ (.A(_3174_),
    .B(_1594_),
    .CON(_0749_),
    .SN(_3544_));
 HAxp5_ASAP7_75t_R _6796_ (.A(_3171_),
    .B(_3545_),
    .CON(_0750_),
    .SN(_0055_));
 HAxp5_ASAP7_75t_R _6797_ (.A(_1207_),
    .B(_3546_),
    .CON(_0107_),
    .SN(_0057_));
 HAxp5_ASAP7_75t_R _6798_ (.A(_1314_),
    .B(_3547_),
    .CON(_0105_),
    .SN(_0751_));
 HAxp5_ASAP7_75t_R _6799_ (.A(_1336_),
    .B(_3548_),
    .CON(_0106_),
    .SN(_0062_));
 HAxp5_ASAP7_75t_R _6800_ (.A(_1388_),
    .B(_3549_),
    .CON(_0101_),
    .SN(_0752_));
 HAxp5_ASAP7_75t_R _6801_ (.A(_3244_),
    .B(_3550_),
    .CON(_0102_),
    .SN(_0069_));
 HAxp5_ASAP7_75t_R _6802_ (.A(_3436_),
    .B(_3551_),
    .CON(_0103_),
    .SN(_0753_));
 HAxp5_ASAP7_75t_R _6803_ (.A(_3442_),
    .B(_3552_),
    .CON(_0104_),
    .SN(_0072_));
 HAxp5_ASAP7_75t_R _6804_ (.A(_3553_),
    .B(_3554_),
    .CON(_0754_),
    .SN(_0080_));
 HAxp5_ASAP7_75t_R _6805_ (.A(_3154_),
    .B(_3555_),
    .CON(_0096_),
    .SN(_0083_));
 HAxp5_ASAP7_75t_R _6806_ (.A(_1348_),
    .B(_3556_),
    .CON(_0097_),
    .SN(_0755_));
 HAxp5_ASAP7_75t_R _6807_ (.A(_3239_),
    .B(_3557_),
    .CON(_0098_),
    .SN(_0084_));
 HAxp5_ASAP7_75t_R _6808_ (.A(_3191_),
    .B(_3558_),
    .CON(_0099_),
    .SN(_0756_));
 HAxp5_ASAP7_75t_R _6809_ (.A(_3468_),
    .B(_3559_),
    .CON(_0100_),
    .SN(_0087_));
 HAxp5_ASAP7_75t_R _6810_ (.A(_3560_),
    .B(_3561_),
    .CON(_0757_),
    .SN(_0088_));
 HAxp5_ASAP7_75t_R _6811_ (.A(_3562_),
    .B(_3563_),
    .CON(_0758_),
    .SN(_0089_));
 HAxp5_ASAP7_75t_R _6812_ (.A(_3564_),
    .B(_3565_),
    .CON(_0759_),
    .SN(_0090_));
 HAxp5_ASAP7_75t_R _6813_ (.A(_3566_),
    .B(_3567_),
    .CON(_0760_),
    .SN(_0091_));
 HAxp5_ASAP7_75t_R _6814_ (.A(_3568_),
    .B(_3569_),
    .CON(_0761_),
    .SN(_0092_));
 HAxp5_ASAP7_75t_R _6815_ (.A(_3570_),
    .B(_3571_),
    .CON(_0762_),
    .SN(_0093_));
 HAxp5_ASAP7_75t_R _6816_ (.A(_3572_),
    .B(_3573_),
    .CON(_0763_),
    .SN(_0094_));
 HAxp5_ASAP7_75t_R _6817_ (.A(_3574_),
    .B(_3575_),
    .CON(_0764_),
    .SN(_0095_));
 HAxp5_ASAP7_75t_R _6818_ (.A(\__st_0[3] ),
    .B(_3576_),
    .CON(_0109_),
    .SN(_0765_));
 HAxp5_ASAP7_75t_R _6819_ (.A(_1677_),
    .B(_1877_),
    .CON(_0108_),
    .SN(_0110_));
 HAxp5_ASAP7_75t_R _6820_ (.A(\__st_0[2] ),
    .B(_3579_),
    .CON(_0111_),
    .SN(_0112_));
 HAxp5_ASAP7_75t_R _6821_ (.A(\__st_0[6] ),
    .B(_3580_),
    .CON(_0766_),
    .SN(_0113_));
 HAxp5_ASAP7_75t_R _6822_ (.A(\__st_0[4] ),
    .B(_3581_),
    .CON(_0114_),
    .SN(_0115_));
 HAxp5_ASAP7_75t_R _6823_ (.A(_3409_),
    .B(_1207_),
    .CON(_0767_),
    .SN(_0117_));
 HAxp5_ASAP7_75t_R _6824_ (.A(_3217_),
    .B(_1882_),
    .CON(_0768_),
    .SN(_0118_));
 HAxp5_ASAP7_75t_R _6825_ (.A(_3233_),
    .B(_3583_),
    .CON(_0769_),
    .SN(_0119_));
 HAxp5_ASAP7_75t_R _6826_ (.A(_3584_),
    .B(_3585_),
    .CON(_3646_),
    .SN(_0120_));
 HAxp5_ASAP7_75t_R _6827_ (.A(_3154_),
    .B(_3191_),
    .CON(_0121_),
    .SN(_0770_));
 HAxp5_ASAP7_75t_R _6828_ (.A(_1348_),
    .B(_3468_),
    .CON(_0122_),
    .SN(_0123_));
 HAxp5_ASAP7_75t_R _6829_ (.A(_3239_),
    .B(_1388_),
    .CON(_0124_),
    .SN(_0771_));
 HAxp5_ASAP7_75t_R _6830_ (.A(_3191_),
    .B(_3244_),
    .CON(_0125_),
    .SN(_0126_));
 HAxp5_ASAP7_75t_R _6831_ (.A(_3436_),
    .B(_3468_),
    .CON(_0127_),
    .SN(_0772_));
 HAxp5_ASAP7_75t_R _6832_ (.A(_3442_),
    .B(_1388_),
    .CON(_0128_),
    .SN(_0129_));
 HAxp5_ASAP7_75t_R _6833_ (.A(_1314_),
    .B(_3244_),
    .CON(_0130_),
    .SN(_0773_));
 HAxp5_ASAP7_75t_R _6834_ (.A(_3436_),
    .B(_1336_),
    .CON(_0131_),
    .SN(_0132_));
 HAxp5_ASAP7_75t_R _6835_ (.A(_1207_),
    .B(_3442_),
    .CON(_0133_),
    .SN(_0774_));
 HAxp5_ASAP7_75t_R _6836_ (.A(_3233_),
    .B(_1314_),
    .CON(_0134_),
    .SN(_0135_));
 HAxp5_ASAP7_75t_R _6837_ (.A(_3154_),
    .B(_3586_),
    .CON(_0136_),
    .SN(_0137_));
 HAxp5_ASAP7_75t_R _6838_ (.A(_3154_),
    .B(_3587_),
    .CON(_0138_),
    .SN(_0775_));
 HAxp5_ASAP7_75t_R _6839_ (.A(_3239_),
    .B(_3588_),
    .CON(_0776_),
    .SN(_0139_));
 HAxp5_ASAP7_75t_R _6840_ (.A(_1348_),
    .B(_3221_),
    .CON(_0140_),
    .SN(_0141_));
 HAxp5_ASAP7_75t_R _6841_ (.A(_3239_),
    .B(_3589_),
    .CON(_0142_),
    .SN(_0777_));
 HAxp5_ASAP7_75t_R _6842_ (.A(_3191_),
    .B(_1897_),
    .CON(_0143_),
    .SN(_0144_));
 HAxp5_ASAP7_75t_R _6843_ (.A(_3468_),
    .B(_3591_),
    .CON(_0145_),
    .SN(_0778_));
 HAxp5_ASAP7_75t_R _6844_ (.A(_1388_),
    .B(_1899_),
    .CON(_0146_),
    .SN(_0147_));
 HAxp5_ASAP7_75t_R _6845_ (.A(_3244_),
    .B(_3593_),
    .CON(_0148_),
    .SN(_0779_));
 HAxp5_ASAP7_75t_R _6846_ (.A(_3436_),
    .B(_1901_),
    .CON(_0149_),
    .SN(_0150_));
 HAxp5_ASAP7_75t_R _6847_ (.A(_3442_),
    .B(_3595_),
    .CON(_0151_),
    .SN(_0780_));
 HAxp5_ASAP7_75t_R _6848_ (.A(_1314_),
    .B(_1904_),
    .CON(_0152_),
    .SN(_0153_));
 HAxp5_ASAP7_75t_R _6849_ (.A(_1336_),
    .B(_2125_),
    .CON(_0154_),
    .SN(_0781_));
 HAxp5_ASAP7_75t_R _6850_ (.A(_1207_),
    .B(_1906_),
    .CON(_0155_),
    .SN(_0156_));
 HAxp5_ASAP7_75t_R _6851_ (.A(_3599_),
    .B(_3600_),
    .CON(_0782_),
    .SN(_0158_));
 HAxp5_ASAP7_75t_R _6852_ (.A(_3154_),
    .B(_1932_),
    .CON(_0161_),
    .SN(_0162_));
 HAxp5_ASAP7_75t_R _6853_ (.A(_1348_),
    .B(_3601_),
    .CON(_0163_),
    .SN(_0783_));
 HAxp5_ASAP7_75t_R _6854_ (.A(_3239_),
    .B(_3240_),
    .CON(_0164_),
    .SN(_0165_));
 HAxp5_ASAP7_75t_R _6855_ (.A(_3191_),
    .B(_1980_),
    .CON(_0166_),
    .SN(_0784_));
 HAxp5_ASAP7_75t_R _6856_ (.A(_3468_),
    .B(_3603_),
    .CON(_0167_),
    .SN(_0168_));
 HAxp5_ASAP7_75t_R _6857_ (.A(_1388_),
    .B(_1986_),
    .CON(_0169_),
    .SN(_0785_));
 HAxp5_ASAP7_75t_R _6858_ (.A(_3244_),
    .B(_3245_),
    .CON(_0170_),
    .SN(_0171_));
 HAxp5_ASAP7_75t_R _6859_ (.A(_3436_),
    .B(_3605_),
    .CON(_0172_),
    .SN(_0786_));
 HAxp5_ASAP7_75t_R _6860_ (.A(_3442_),
    .B(_3606_),
    .CON(_0173_),
    .SN(_0174_));
 HAxp5_ASAP7_75t_R _6861_ (.A(_1314_),
    .B(_3607_),
    .CON(_0175_),
    .SN(_0787_));
 HAxp5_ASAP7_75t_R _6862_ (.A(_1336_),
    .B(_3608_),
    .CON(_0176_),
    .SN(_0177_));
 HAxp5_ASAP7_75t_R _6863_ (.A(_3609_),
    .B(_3610_),
    .CON(_0179_),
    .SN(_0180_));
 HAxp5_ASAP7_75t_R _6864_ (.A(_3611_),
    .B(_3612_),
    .CON(_0788_),
    .SN(_0789_));
 HAxp5_ASAP7_75t_R _6865_ (.A(\__st_1[29] ),
    .B(_3260_),
    .CON(_0790_),
    .SN(_0189_));
 HAxp5_ASAP7_75t_R _6866_ (.A(\__st_1[28] ),
    .B(_3260_),
    .CON(_0190_),
    .SN(_0191_));
 HAxp5_ASAP7_75t_R _6867_ (.A(\__st_1[27] ),
    .B(_3260_),
    .CON(_0791_),
    .SN(_0192_));
 HAxp5_ASAP7_75t_R _6868_ (.A(\__st_1[26] ),
    .B(_3260_),
    .CON(_0193_),
    .SN(_0194_));
 HAxp5_ASAP7_75t_R _6869_ (.A(\__st_1[25] ),
    .B(_3260_),
    .CON(_0792_),
    .SN(_0195_));
 HAxp5_ASAP7_75t_R _6870_ (.A(\__st_1[24] ),
    .B(_3260_),
    .CON(_0196_),
    .SN(_0197_));
 HAxp5_ASAP7_75t_R _6871_ (.A(\__st_1[23] ),
    .B(_3260_),
    .CON(_0198_),
    .SN(_0793_));
 HAxp5_ASAP7_75t_R _6872_ (.A(\__st_1[22] ),
    .B(_3260_),
    .CON(_0199_),
    .SN(_0200_));
 HAxp5_ASAP7_75t_R _6873_ (.A(\__st_1[21] ),
    .B(_3260_),
    .CON(_0794_),
    .SN(_0201_));
 HAxp5_ASAP7_75t_R _6874_ (.A(\__st_1[20] ),
    .B(_3260_),
    .CON(_0202_),
    .SN(_0203_));
 HAxp5_ASAP7_75t_R _6875_ (.A(\__st_1[19] ),
    .B(_3260_),
    .CON(_0204_),
    .SN(_0795_));
 HAxp5_ASAP7_75t_R _6876_ (.A(\__st_1[18] ),
    .B(_3260_),
    .CON(_0205_),
    .SN(_0206_));
 HAxp5_ASAP7_75t_R _6877_ (.A(\__st_1[17] ),
    .B(_3613_),
    .CON(_0207_),
    .SN(_0796_));
 HAxp5_ASAP7_75t_R _6878_ (.A(_3614_),
    .B(_3615_),
    .CON(_0797_),
    .SN(_0208_));
 HAxp5_ASAP7_75t_R _6879_ (.A(\__st_1[16] ),
    .B(_3616_),
    .CON(_0209_),
    .SN(_0210_));
 HAxp5_ASAP7_75t_R _6880_ (.A(\__st_1[15] ),
    .B(_3617_),
    .CON(_0212_),
    .SN(_0798_));
 HAxp5_ASAP7_75t_R _6881_ (.A(_2055_),
    .B(_3619_),
    .CON(_0211_),
    .SN(_0213_));
 HAxp5_ASAP7_75t_R _6882_ (.A(\__st_1[14] ),
    .B(_3283_),
    .CON(_0214_),
    .SN(_0215_));
 HAxp5_ASAP7_75t_R _6883_ (.A(\__st_1[13] ),
    .B(_3620_),
    .CON(_0216_),
    .SN(_0799_));
 HAxp5_ASAP7_75t_R _6884_ (.A(_3621_),
    .B(_3622_),
    .CON(_0800_),
    .SN(_0217_));
 HAxp5_ASAP7_75t_R _6885_ (.A(\__st_1[12] ),
    .B(_3623_),
    .CON(_0218_),
    .SN(_0219_));
 HAxp5_ASAP7_75t_R _6886_ (.A(\__st_1[11] ),
    .B(_3624_),
    .CON(_0220_),
    .SN(_0801_));
 HAxp5_ASAP7_75t_R _6887_ (.A(_3625_),
    .B(_3626_),
    .CON(_0802_),
    .SN(_0221_));
 HAxp5_ASAP7_75t_R _6888_ (.A(\__st_1[10] ),
    .B(_3627_),
    .CON(_0222_),
    .SN(_0223_));
 HAxp5_ASAP7_75t_R _6889_ (.A(\__st_1[9] ),
    .B(_3628_),
    .CON(_0224_),
    .SN(_0803_));
 HAxp5_ASAP7_75t_R _6890_ (.A(_3629_),
    .B(_3630_),
    .CON(_0804_),
    .SN(_0225_));
 HAxp5_ASAP7_75t_R _6891_ (.A(\__st_1[8] ),
    .B(_3631_),
    .CON(_0226_),
    .SN(_0227_));
 HAxp5_ASAP7_75t_R _6892_ (.A(\__st_1[7] ),
    .B(_3632_),
    .CON(_0228_),
    .SN(_0805_));
 HAxp5_ASAP7_75t_R _6893_ (.A(_3633_),
    .B(_3634_),
    .CON(_0806_),
    .SN(_0229_));
 HAxp5_ASAP7_75t_R _6894_ (.A(\__st_1[6] ),
    .B(_3635_),
    .CON(_0230_),
    .SN(_0231_));
 HAxp5_ASAP7_75t_R _6895_ (.A(\__st_1[5] ),
    .B(_3636_),
    .CON(_0232_),
    .SN(_0807_));
 HAxp5_ASAP7_75t_R _6896_ (.A(_3637_),
    .B(_3638_),
    .CON(_0808_),
    .SN(_0233_));
 HAxp5_ASAP7_75t_R _6897_ (.A(\__st_1[4] ),
    .B(_3639_),
    .CON(_0234_),
    .SN(_0235_));
 HAxp5_ASAP7_75t_R _6898_ (.A(\__st_1[3] ),
    .B(_3640_),
    .CON(_0236_),
    .SN(_0809_));
 HAxp5_ASAP7_75t_R _6899_ (.A(_3641_),
    .B(_3642_),
    .CON(_0810_),
    .SN(_0237_));
 HAxp5_ASAP7_75t_R _6900_ (.A(\__st_1[2] ),
    .B(_3643_),
    .CON(_0238_),
    .SN(_0239_));
 HAxp5_ASAP7_75t_R _6901_ (.A(_3644_),
    .B(_3645_),
    .CON(_0811_),
    .SN(_0240_));
 HAxp5_ASAP7_75t_R _6902_ (.A(\__st_2[0] ),
    .B(net229),
    .CON(_0812_),
    .SN(_0813_));
 HAxp5_ASAP7_75t_R _6903_ (.A(\__st_2[13] ),
    .B(net229),
    .CON(_0244_),
    .SN(_0814_));
 HAxp5_ASAP7_75t_R _6904_ (.A(\__st_2[12] ),
    .B(net229),
    .CON(_0245_),
    .SN(_0246_));
 HAxp5_ASAP7_75t_R _6905_ (.A(\__st_2[11] ),
    .B(net229),
    .CON(_0247_),
    .SN(_0815_));
 HAxp5_ASAP7_75t_R _6906_ (.A(\__st_2[10] ),
    .B(net229),
    .CON(_0248_),
    .SN(_0249_));
 HAxp5_ASAP7_75t_R _6907_ (.A(\__st_2[9] ),
    .B(net229),
    .CON(_0250_),
    .SN(_0251_));
 HAxp5_ASAP7_75t_R _6908_ (.A(\__st_2[8] ),
    .B(net229),
    .CON(_0252_),
    .SN(_0253_));
 HAxp5_ASAP7_75t_R _6909_ (.A(\__st_2[7] ),
    .B(net229),
    .CON(_0254_),
    .SN(_0255_));
 HAxp5_ASAP7_75t_R _6910_ (.A(\__st_2[3] ),
    .B(_3576_),
    .CON(_0256_),
    .SN(_0816_));
 HAxp5_ASAP7_75t_R _6911_ (.A(\__st_2[2] ),
    .B(_3579_),
    .CON(_0257_),
    .SN(_0258_));
 HAxp5_ASAP7_75t_R _6912_ (.A(\__st_2[6] ),
    .B(_3648_),
    .CON(_0817_),
    .SN(_0260_));
 HAxp5_ASAP7_75t_R _6913_ (.A(\__st_2[4] ),
    .B(_3649_),
    .CON(_0261_),
    .SN(_0262_));
 HAxp5_ASAP7_75t_R _6914_ (.A(_3650_),
    .B(_3651_),
    .CON(_0818_),
    .SN(_0265_));
 HAxp5_ASAP7_75t_R _6915_ (.A(_3652_),
    .B(_3653_),
    .CON(_0819_),
    .SN(_0820_));
 HAxp5_ASAP7_75t_R _6916_ (.A(_3654_),
    .B(_3655_),
    .CON(_0821_),
    .SN(_0266_));
 HAxp5_ASAP7_75t_R _6917_ (.A(_3656_),
    .B(_2209_),
    .CON(_0822_),
    .SN(_0267_));
 HAxp5_ASAP7_75t_R _6918_ (.A(_3337_),
    .B(_2261_),
    .CON(_0268_),
    .SN(_0823_));
 HAxp5_ASAP7_75t_R _6919_ (.A(_2220_),
    .B(_2271_),
    .CON(_0269_),
    .SN(_0270_));
 HAxp5_ASAP7_75t_R _6920_ (.A(_2240_),
    .B(_2290_),
    .CON(_0271_),
    .SN(_0824_));
 HAxp5_ASAP7_75t_R _6921_ (.A(_2261_),
    .B(_2315_),
    .CON(_0272_),
    .SN(_0273_));
 HAxp5_ASAP7_75t_R _6922_ (.A(_2271_),
    .B(_2333_),
    .CON(_0274_),
    .SN(_0825_));
 HAxp5_ASAP7_75t_R _6923_ (.A(_2290_),
    .B(_3348_),
    .CON(_0275_),
    .SN(_0276_));
 HAxp5_ASAP7_75t_R _6924_ (.A(_2315_),
    .B(_3325_),
    .CON(_0277_),
    .SN(_0826_));
 HAxp5_ASAP7_75t_R _6925_ (.A(_2333_),
    .B(_2417_),
    .CON(_0278_),
    .SN(_0279_));
 HAxp5_ASAP7_75t_R _6926_ (.A(_3348_),
    .B(_2436_),
    .CON(_0280_),
    .SN(_0827_));
 HAxp5_ASAP7_75t_R _6927_ (.A(_3325_),
    .B(_2459_),
    .CON(_0281_),
    .SN(_0282_));
 HAxp5_ASAP7_75t_R _6928_ (.A(_3337_),
    .B(_3659_),
    .CON(_0283_),
    .SN(_0284_));
 HAxp5_ASAP7_75t_R _6929_ (.A(_3337_),
    .B(_3660_),
    .CON(_0286_),
    .SN(_0828_));
 HAxp5_ASAP7_75t_R _6930_ (.A(_2240_),
    .B(_3661_),
    .CON(_0829_),
    .SN(_0287_));
 HAxp5_ASAP7_75t_R _6931_ (.A(_2220_),
    .B(_3316_),
    .CON(_0288_),
    .SN(_0289_));
 HAxp5_ASAP7_75t_R _6932_ (.A(_2240_),
    .B(_3662_),
    .CON(_0830_),
    .SN(_0831_));
 HAxp5_ASAP7_75t_R _6933_ (.A(_2261_),
    .B(_3318_),
    .CON(_0290_),
    .SN(_0291_));
 HAxp5_ASAP7_75t_R _6934_ (.A(_2271_),
    .B(_2595_),
    .CON(_0292_),
    .SN(_0832_));
 HAxp5_ASAP7_75t_R _6935_ (.A(_2290_),
    .B(_2551_),
    .CON(_0293_),
    .SN(_0294_));
 HAxp5_ASAP7_75t_R _6936_ (.A(_2315_),
    .B(_2583_),
    .CON(_0295_),
    .SN(_0833_));
 HAxp5_ASAP7_75t_R _6937_ (.A(_2333_),
    .B(_2558_),
    .CON(_0296_),
    .SN(_0297_));
 HAxp5_ASAP7_75t_R _6938_ (.A(_3348_),
    .B(_3665_),
    .CON(_0299_),
    .SN(_0834_));
 HAxp5_ASAP7_75t_R _6939_ (.A(_3325_),
    .B(_3326_),
    .CON(_0301_),
    .SN(_0302_));
 HAxp5_ASAP7_75t_R _6940_ (.A(_2417_),
    .B(_3666_),
    .CON(_0303_),
    .SN(_0835_));
 HAxp5_ASAP7_75t_R _6941_ (.A(_2436_),
    .B(_3668_),
    .CON(_0304_),
    .SN(_0305_));
 HAxp5_ASAP7_75t_R _6942_ (.A(_2436_),
    .B(_3669_),
    .CON(_3312_),
    .SN(_0306_));
 HAxp5_ASAP7_75t_R _6943_ (.A(_3670_),
    .B(_3671_),
    .CON(_0836_),
    .SN(_0307_));
 HAxp5_ASAP7_75t_R _6944_ (.A(_3337_),
    .B(_3338_),
    .CON(_0308_),
    .SN(_0309_));
 HAxp5_ASAP7_75t_R _6945_ (.A(_2220_),
    .B(_3672_),
    .CON(_0837_),
    .SN(_0838_));
 HAxp5_ASAP7_75t_R _6946_ (.A(_2240_),
    .B(_2547_),
    .CON(_0312_),
    .SN(_0313_));
 HAxp5_ASAP7_75t_R _6947_ (.A(_2261_),
    .B(_3673_),
    .CON(_0315_),
    .SN(_0839_));
 HAxp5_ASAP7_75t_R _6948_ (.A(_2271_),
    .B(_2553_),
    .CON(_0317_),
    .SN(_0318_));
 HAxp5_ASAP7_75t_R _6949_ (.A(_2290_),
    .B(_3674_),
    .CON(_0320_),
    .SN(_0840_));
 HAxp5_ASAP7_75t_R _6950_ (.A(_2315_),
    .B(_3346_),
    .CON(_0322_),
    .SN(_0323_));
 HAxp5_ASAP7_75t_R _6951_ (.A(_2333_),
    .B(_3675_),
    .CON(_0325_),
    .SN(_0841_));
 HAxp5_ASAP7_75t_R _6952_ (.A(_3348_),
    .B(_2566_),
    .CON(_0327_),
    .SN(_0328_));
 HAxp5_ASAP7_75t_R _6953_ (.A(_3325_),
    .B(_3676_),
    .CON(_0329_),
    .SN(_0842_));
 HAxp5_ASAP7_75t_R _6954_ (.A(_2417_),
    .B(_3678_),
    .CON(_0330_),
    .SN(_0331_));
 HAxp5_ASAP7_75t_R _6955_ (.A(_3658_),
    .B(_3679_),
    .CON(_3332_),
    .SN(_0332_));
 HAxp5_ASAP7_75t_R _6956_ (.A(_3680_),
    .B(_3681_),
    .CON(_0843_),
    .SN(_0844_));
 HAxp5_ASAP7_75t_R _6957_ (.A(_2459_),
    .B(_3682_),
    .CON(_0845_),
    .SN(_0342_));
 HAxp5_ASAP7_75t_R _6958_ (.A(net27),
    .B(_3683_),
    .CON(_0407_),
    .SN(_0344_));
 HAxp5_ASAP7_75t_R _6959_ (.A(_3684_),
    .B(_3685_),
    .CON(_0846_),
    .SN(_0345_));
 HAxp5_ASAP7_75t_R _6960_ (.A(net26),
    .B(_3686_),
    .CON(_0346_),
    .SN(_0347_));
 HAxp5_ASAP7_75t_R _6961_ (.A(net25),
    .B(_3687_),
    .CON(_0847_),
    .SN(_0848_));
 HAxp5_ASAP7_75t_R _6962_ (.A(_3688_),
    .B(_3689_),
    .CON(_0849_),
    .SN(_0348_));
 HAxp5_ASAP7_75t_R _6963_ (.A(net24),
    .B(_3690_),
    .CON(_0349_),
    .SN(_0351_));
 HAxp5_ASAP7_75t_R _6964_ (.A(net23),
    .B(_3691_),
    .CON(_0850_),
    .SN(_0851_));
 HAxp5_ASAP7_75t_R _6965_ (.A(_3692_),
    .B(_3693_),
    .CON(_0852_),
    .SN(_0353_));
 HAxp5_ASAP7_75t_R _6966_ (.A(net22),
    .B(_3694_),
    .CON(_0354_),
    .SN(_0355_));
 HAxp5_ASAP7_75t_R _6967_ (.A(net36),
    .B(_3695_),
    .CON(_0357_),
    .SN(_0853_));
 HAxp5_ASAP7_75t_R _6968_ (.A(_3696_),
    .B(_3697_),
    .CON(_0854_),
    .SN(_0358_));
 HAxp5_ASAP7_75t_R _6969_ (.A(net35),
    .B(_3698_),
    .CON(_0359_),
    .SN(_0360_));
 HAxp5_ASAP7_75t_R _6970_ (.A(net34),
    .B(_3699_),
    .CON(_0361_),
    .SN(_0855_));
 HAxp5_ASAP7_75t_R _6971_ (.A(_3700_),
    .B(_3701_),
    .CON(_0856_),
    .SN(_0362_));
 HAxp5_ASAP7_75t_R _6972_ (.A(net33),
    .B(_3702_),
    .CON(_0363_),
    .SN(_0364_));
 HAxp5_ASAP7_75t_R _6973_ (.A(net32),
    .B(_3703_),
    .CON(_0365_),
    .SN(_0857_));
 HAxp5_ASAP7_75t_R _6974_ (.A(_3704_),
    .B(_2667_),
    .CON(_0858_),
    .SN(_0367_));
 HAxp5_ASAP7_75t_R _6975_ (.A(net31),
    .B(_3706_),
    .CON(_0368_),
    .SN(_0369_));
 HAxp5_ASAP7_75t_R _6976_ (.A(net30),
    .B(_3707_),
    .CON(_0370_),
    .SN(_0859_));
 HAxp5_ASAP7_75t_R _6977_ (.A(_3708_),
    .B(_3709_),
    .CON(_0860_),
    .SN(_0371_));
 HAxp5_ASAP7_75t_R _6978_ (.A(net29),
    .B(_3710_),
    .CON(_0372_),
    .SN(_0374_));
 HAxp5_ASAP7_75t_R _6979_ (.A(_3711_),
    .B(_3712_),
    .CON(_0343_),
    .SN(_0375_));
 HAxp5_ASAP7_75t_R _6980_ (.A(_3713_),
    .B(_3714_),
    .CON(_0378_),
    .SN(_0379_));
 HAxp5_ASAP7_75t_R _6981_ (.A(\__st_3[29] ),
    .B(_3365_),
    .CON(_0861_),
    .SN(_0381_));
 HAxp5_ASAP7_75t_R _6982_ (.A(\__st_3[28] ),
    .B(_3365_),
    .CON(_0382_),
    .SN(_0383_));
 HAxp5_ASAP7_75t_R _6983_ (.A(\__st_3[27] ),
    .B(_3365_),
    .CON(_0862_),
    .SN(_0384_));
 HAxp5_ASAP7_75t_R _6984_ (.A(\__st_3[26] ),
    .B(_3365_),
    .CON(_0385_),
    .SN(_0386_));
 HAxp5_ASAP7_75t_R _6985_ (.A(\__st_3[25] ),
    .B(_3365_),
    .CON(_0863_),
    .SN(_0387_));
 HAxp5_ASAP7_75t_R _6986_ (.A(\__st_3[24] ),
    .B(_3365_),
    .CON(_0388_),
    .SN(_0390_));
 HAxp5_ASAP7_75t_R _6987_ (.A(\__st_3[23] ),
    .B(_3365_),
    .CON(_0391_),
    .SN(_0864_));
 HAxp5_ASAP7_75t_R _6988_ (.A(\__st_3[22] ),
    .B(_3365_),
    .CON(_0393_),
    .SN(_0394_));
 HAxp5_ASAP7_75t_R _6989_ (.A(\__st_3[21] ),
    .B(_3365_),
    .CON(_0395_),
    .SN(_0865_));
 HAxp5_ASAP7_75t_R _6990_ (.A(\__st_3[20] ),
    .B(_3365_),
    .CON(_0396_),
    .SN(_0398_));
 HAxp5_ASAP7_75t_R _6991_ (.A(\__st_3[19] ),
    .B(_3365_),
    .CON(_0399_),
    .SN(_0866_));
 HAxp5_ASAP7_75t_R _6992_ (.A(\__st_3[18] ),
    .B(_3365_),
    .CON(_0400_),
    .SN(_0401_));
 HAxp5_ASAP7_75t_R _6993_ (.A(\__st_3[17] ),
    .B(_3715_),
    .CON(_0402_),
    .SN(_0403_));
 HAxp5_ASAP7_75t_R _6994_ (.A(_3716_),
    .B(_3717_),
    .CON(_0867_),
    .SN(_0404_));
 HAxp5_ASAP7_75t_R _6995_ (.A(\__st_3[16] ),
    .B(_3371_),
    .CON(_0405_),
    .SN(_0406_));
 HAxp5_ASAP7_75t_R _6996_ (.A(_3718_),
    .B(_3719_),
    .CON(_3720_),
    .SN(_0414_));
 DFFLQNx2_ASAP7_75t_R _6997_ (.QN(_3584_),
    .CLK(net161),
    .D(_0869_));
 DFFLQNx2_ASAP7_75t_R _6998_ (.QN(_3123_),
    .CLK(net160),
    .D(_0870_));
 DFFLQNx2_ASAP7_75t_R _6999_ (.QN(_3126_),
    .CLK(net159),
    .D(_0871_));
 DFFLQNx2_ASAP7_75t_R _7000_ (.QN(_3426_),
    .CLK(net158),
    .D(_0872_));
 DFFLQNx2_ASAP7_75t_R _7001_ (.QN(_3272_),
    .CLK(net157),
    .D(_0873_));
 DFFLQNx2_ASAP7_75t_R _7002_ (.QN(_3425_),
    .CLK(net156),
    .D(_0874_));
 DFFLQNx2_ASAP7_75t_R _7003_ (.QN(_3127_),
    .CLK(net155),
    .D(_0875_));
 DFFLQNx2_ASAP7_75t_R _7004_ (.QN(_3424_),
    .CLK(net154),
    .D(_0876_));
 DFFLQNx2_ASAP7_75t_R _7005_ (.QN(_3137_),
    .CLK(net153),
    .D(_0877_));
 DFFLQNx2_ASAP7_75t_R _7006_ (.QN(_3423_),
    .CLK(net152),
    .D(_0878_));
 DFFLQNx2_ASAP7_75t_R _7007_ (.QN(_3135_),
    .CLK(net151),
    .D(_0879_));
 DFFLQNx2_ASAP7_75t_R _7008_ (.QN(_3422_),
    .CLK(net150),
    .D(_0880_));
 DFFLQNx2_ASAP7_75t_R _7009_ (.QN(_3133_),
    .CLK(net149),
    .D(_0881_));
 DFFLQNx2_ASAP7_75t_R _7010_ (.QN(_3421_),
    .CLK(net148),
    .D(_0882_));
 DFFLQNx2_ASAP7_75t_R _7011_ (.QN(_3131_),
    .CLK(net147),
    .D(_0883_));
 DFFLQNx2_ASAP7_75t_R _7012_ (.QN(_3420_),
    .CLK(net146),
    .D(_0884_));
 DFFLQNx2_ASAP7_75t_R _7013_ (.QN(_3265_),
    .CLK(net145),
    .D(_0885_));
 DFFLQNx2_ASAP7_75t_R _7014_ (.QN(_3419_),
    .CLK(net144),
    .D(_0886_));
 DFFLQNx2_ASAP7_75t_R _7015_ (.QN(_3418_),
    .CLK(net143),
    .D(_0887_));
 DFFLQNx2_ASAP7_75t_R _7016_ (.QN(_3417_),
    .CLK(net142),
    .D(_0888_));
 DFFLQNx2_ASAP7_75t_R _7017_ (.QN(_3262_),
    .CLK(net141),
    .D(_0889_));
 DFFLQNx2_ASAP7_75t_R _7018_ (.QN(_3416_),
    .CLK(net140),
    .D(_0890_));
 DFFLQNx2_ASAP7_75t_R _7019_ (.QN(_3415_),
    .CLK(net139),
    .D(_0891_));
 DFFLQNx2_ASAP7_75t_R _7020_ (.QN(_3414_),
    .CLK(net138),
    .D(_0892_));
 DFFLQNx2_ASAP7_75t_R _7021_ (.QN(_3258_),
    .CLK(net137),
    .D(_0893_));
 DFFLQNx2_ASAP7_75t_R _7022_ (.QN(_3413_),
    .CLK(net136),
    .D(_0894_));
 DFFLQNx2_ASAP7_75t_R _7023_ (.QN(_3143_),
    .CLK(net135),
    .D(_0895_));
 DFFLQNx2_ASAP7_75t_R _7024_ (.QN(_3412_),
    .CLK(net134),
    .D(_0896_));
 DFFLQNx2_ASAP7_75t_R _7025_ (.QN(_3141_),
    .CLK(net133),
    .D(_0897_));
 DFFLQNx2_ASAP7_75t_R _7026_ (.QN(_3411_),
    .CLK(net132),
    .D(_0898_));
 DFFLQNx2_ASAP7_75t_R _7027_ (.QN(_3139_),
    .CLK(net131),
    .D(_0899_));
 DFFLQNx2_ASAP7_75t_R _7028_ (.QN(_0567_),
    .CLK(net130),
    .D(_0900_));
 DFFLQNx2_ASAP7_75t_R _7029_ (.QN(_0566_),
    .CLK(net129),
    .D(_0901_));
 DFFLQNx2_ASAP7_75t_R _7030_ (.QN(_0565_),
    .CLK(net128),
    .D(_0902_));
 DFFLQNx2_ASAP7_75t_R _7031_ (.QN(_3292_),
    .CLK(net127),
    .D(_0903_));
 DFFLQNx2_ASAP7_75t_R _7032_ (.QN(_0564_),
    .CLK(net126),
    .D(_0904_));
 DFFLQNx2_ASAP7_75t_R _7033_ (.QN(_0563_),
    .CLK(net125),
    .D(_0905_));
 DFFLQNx2_ASAP7_75t_R _7034_ (.QN(_0562_),
    .CLK(net124),
    .D(_0906_));
 DFFLQNx2_ASAP7_75t_R _7035_ (.QN(_0259_),
    .CLK(net123),
    .D(_0907_));
 DFFLQNx2_ASAP7_75t_R _7036_ (.QN(_0561_),
    .CLK(net122),
    .D(_0908_));
 DFFLQNx2_ASAP7_75t_R _7037_ (.QN(_0560_),
    .CLK(net121),
    .D(_0909_));
 DFFLQNx2_ASAP7_75t_R _7038_ (.QN(_0559_),
    .CLK(net120),
    .D(_0910_));
 DFFLQNx2_ASAP7_75t_R _7039_ (.QN(_3289_),
    .CLK(net119),
    .D(_0911_));
 DFFLQNx2_ASAP7_75t_R _7040_ (.QN(_0558_),
    .CLK(net118),
    .D(_0912_));
 DFFLQNx2_ASAP7_75t_R _7041_ (.QN(_3287_),
    .CLK(net117),
    .D(_0913_));
 DFFLQNx2_ASAP7_75t_R _7042_ (.QN(_0557_),
    .CLK(net116),
    .D(_0914_));
 DFFLQNx2_ASAP7_75t_R _7043_ (.QN(_3285_),
    .CLK(net115),
    .D(_0915_));
 DFFLQNx2_ASAP7_75t_R _7044_ (.QN(_0556_),
    .CLK(net114),
    .D(_0916_));
 DFFLQNx2_ASAP7_75t_R _7045_ (.QN(_0555_),
    .CLK(net113),
    .D(_0917_));
 DFFLQNx2_ASAP7_75t_R _7046_ (.QN(_3206_),
    .CLK(net112),
    .D(_0918_));
 DFFLQNx2_ASAP7_75t_R _7047_ (.QN(_0554_),
    .CLK(net111),
    .D(_0919_));
 DFFLQNx2_ASAP7_75t_R _7048_ (.QN(_0553_),
    .CLK(net110),
    .D(_0920_));
 DFFLQNx2_ASAP7_75t_R _7049_ (.QN(_0552_),
    .CLK(net109),
    .D(_0921_));
 DFFLQNx2_ASAP7_75t_R _7050_ (.QN(_0551_),
    .CLK(net108),
    .D(_0922_));
 DFFLQNx2_ASAP7_75t_R _7051_ (.QN(_0550_),
    .CLK(net107),
    .D(_0923_));
 DFFLQNx2_ASAP7_75t_R _7052_ (.QN(_0549_),
    .CLK(net106),
    .D(_0924_));
 DFFLQNx2_ASAP7_75t_R _7053_ (.QN(_0548_),
    .CLK(net105),
    .D(_0925_));
 DFFLQNx2_ASAP7_75t_R _7054_ (.QN(_3202_),
    .CLK(net104),
    .D(_0926_));
 DFFLQNx2_ASAP7_75t_R _7055_ (.QN(_0547_),
    .CLK(net103),
    .D(_0927_));
 DFFLQNx2_ASAP7_75t_R _7056_ (.QN(_3200_),
    .CLK(net102),
    .D(_0928_));
 DFFLQNx2_ASAP7_75t_R _7057_ (.QN(_0546_),
    .CLK(net101),
    .D(_0929_));
 DFFLQNx2_ASAP7_75t_R _7058_ (.QN(_3197_),
    .CLK(net100),
    .D(_0930_));
 DFFLQNx2_ASAP7_75t_R _7059_ (.QN(_3718_),
    .CLK(net99),
    .D(_0931_));
 DFFLQNx2_ASAP7_75t_R _7060_ (.QN(_3373_),
    .CLK(net98),
    .D(_0932_));
 DFFLQNx2_ASAP7_75t_R _7061_ (.QN(_3377_),
    .CLK(net97),
    .D(_0933_));
 DFFLQNx2_ASAP7_75t_R _7062_ (.QN(_0545_),
    .CLK(net96),
    .D(_0934_));
 DFFLQNx2_ASAP7_75t_R _7063_ (.QN(_3379_),
    .CLK(net95),
    .D(_0935_));
 DFFLQNx2_ASAP7_75t_R _7064_ (.QN(_0544_),
    .CLK(net94),
    .D(_0936_));
 DFFLQNx2_ASAP7_75t_R _7065_ (.QN(_3382_),
    .CLK(net93),
    .D(_0937_));
 DFFLQNx2_ASAP7_75t_R _7066_ (.QN(_0543_),
    .CLK(net92),
    .D(_0938_));
 DFFLQNx2_ASAP7_75t_R _7067_ (.QN(_3385_),
    .CLK(net91),
    .D(_0939_));
 DFFLQNx2_ASAP7_75t_R _7068_ (.QN(_0542_),
    .CLK(net90),
    .D(_0940_));
 DFFLQNx2_ASAP7_75t_R _7069_ (.QN(_3388_),
    .CLK(net89),
    .D(_0941_));
 DFFLQNx2_ASAP7_75t_R _7070_ (.QN(_0541_),
    .CLK(net88),
    .D(_0942_));
 DFFLQNx2_ASAP7_75t_R _7071_ (.QN(_3391_),
    .CLK(net87),
    .D(_0943_));
 DFFLQNx2_ASAP7_75t_R _7072_ (.QN(_0540_),
    .CLK(net86),
    .D(_0944_));
 DFFLQNx2_ASAP7_75t_R _7073_ (.QN(_3394_),
    .CLK(net85),
    .D(_0945_));
 DFFLQNx2_ASAP7_75t_R _7074_ (.QN(_0539_),
    .CLK(net84),
    .D(_0946_));
 DFFLQNx2_ASAP7_75t_R _7075_ (.QN(_0538_),
    .CLK(net83),
    .D(_0947_));
 DFFLQNx2_ASAP7_75t_R _7076_ (.QN(_0537_),
    .CLK(net82),
    .D(_0948_));
 DFFLQNx2_ASAP7_75t_R _7077_ (.QN(_3369_),
    .CLK(net81),
    .D(_0949_));
 DFFLQNx2_ASAP7_75t_R _7078_ (.QN(_0536_),
    .CLK(net80),
    .D(_0950_));
 DFFLQNx2_ASAP7_75t_R _7079_ (.QN(_3367_),
    .CLK(net79),
    .D(_0951_));
 DFFLQNx2_ASAP7_75t_R _7080_ (.QN(_0535_),
    .CLK(net78),
    .D(_0952_));
 DFFLQNx2_ASAP7_75t_R _7081_ (.QN(_0534_),
    .CLK(net77),
    .D(_0953_));
 DFFLQNx2_ASAP7_75t_R _7082_ (.QN(_0533_),
    .CLK(net76),
    .D(_0954_));
 DFFLQNx2_ASAP7_75t_R _7083_ (.QN(_3363_),
    .CLK(net75),
    .D(_0955_));
 DFFLQNx2_ASAP7_75t_R _7084_ (.QN(_0532_),
    .CLK(net74),
    .D(_0956_));
 DFFLQNx2_ASAP7_75t_R _7085_ (.QN(_3361_),
    .CLK(net73),
    .D(_0957_));
 DFFLQNx2_ASAP7_75t_R _7086_ (.QN(_0531_),
    .CLK(net72),
    .D(_0958_));
 DFFLQNx2_ASAP7_75t_R _7087_ (.QN(_3359_),
    .CLK(net71),
    .D(_0959_));
 DFFLQNx2_ASAP7_75t_R _7088_ (.QN(_0530_),
    .CLK(net70),
    .D(_0960_));
 DFFLQNx2_ASAP7_75t_R _7089_ (.QN(_3356_),
    .CLK(net69),
    .D(_0961_));
 DFFLQNx2_ASAP7_75t_R _7090_ (.QN(_0529_),
    .CLK(net68),
    .D(_0962_));
 DFFLQNx2_ASAP7_75t_R _7091_ (.QN(_3405_),
    .CLK(net67),
    .D(_0963_));
 DFFLQNx2_ASAP7_75t_R _7092_ (.QN(_0528_),
    .CLK(net66),
    .D(_0964_));
 DFFLQNx2_ASAP7_75t_R _7093_ (.QN(_0527_),
    .CLK(net65),
    .D(_0965_));
 DFFLQNx2_ASAP7_75t_R _7094_ (.QN(_0526_),
    .CLK(net64),
    .D(_0966_));
 DFFLQNx2_ASAP7_75t_R _7095_ (.QN(_3129_),
    .CLK(net63),
    .D(_0967_));
 DFFLQNx2_ASAP7_75t_R _7096_ (.QN(_0525_),
    .CLK(net62),
    .D(_0968_));
 DFFLQNx2_ASAP7_75t_R _7097_ (.QN(_0524_),
    .CLK(net61),
    .D(_0969_));
 DFFLQNx2_ASAP7_75t_R _7098_ (.QN(_0523_),
    .CLK(net60),
    .D(_0970_));
 DFFLQNx2_ASAP7_75t_R _7099_ (.QN(_0522_),
    .CLK(net59),
    .D(_0971_));
 DFFLQNx2_ASAP7_75t_R _7100_ (.QN(_0521_),
    .CLK(net58),
    .D(_0972_));
 DFFLQNx2_ASAP7_75t_R _7101_ (.QN(_0520_),
    .CLK(net57),
    .D(_0973_));
 DFFLQNx2_ASAP7_75t_R _7102_ (.QN(_0519_),
    .CLK(net56),
    .D(_0974_));
 DFFLQNx2_ASAP7_75t_R _7103_ (.QN(_0518_),
    .CLK(net55),
    .D(_0975_));
 DFFLQNx2_ASAP7_75t_R _7104_ (.QN(_0517_),
    .CLK(net54),
    .D(_0976_));
 DFFLQNx2_ASAP7_75t_R _7105_ (.QN(_0516_),
    .CLK(net53),
    .D(_0977_));
 DFFLQNx2_ASAP7_75t_R _7106_ (.QN(_3145_),
    .CLK(net52),
    .D(_0978_));
 DFFLQNx2_ASAP7_75t_R _7107_ (.QN(_0427_),
    .CLK(net51),
    .D(_0979_));
 DFFLQNx2_ASAP7_75t_R _7108_ (.QN(_0515_),
    .CLK(net50),
    .D(_0980_));
 TAPCELL_ASAP7_75t_R PHY_15 ();
 TAPCELL_ASAP7_75t_R PHY_14 ();
 TAPCELL_ASAP7_75t_R PHY_13 ();
 TAPCELL_ASAP7_75t_R PHY_12 ();
 TAPCELL_ASAP7_75t_R PHY_11 ();
 TAPCELL_ASAP7_75t_R PHY_10 ();
 TAPCELL_ASAP7_75t_R PHY_9 ();
 TAPCELL_ASAP7_75t_R PHY_8 ();
 TAPCELL_ASAP7_75t_R PHY_7 ();
 TAPCELL_ASAP7_75t_R PHY_6 ();
 TAPCELL_ASAP7_75t_R PHY_5 ();
 TAPCELL_ASAP7_75t_R PHY_4 ();
 TAPCELL_ASAP7_75t_R PHY_3 ();
 TAPCELL_ASAP7_75t_R PHY_2 ();
 TAPCELL_ASAP7_75t_R PHY_1 ();
 TAPCELL_ASAP7_75t_R PHY_0 ();
 BUFx2_ASAP7_75t_R input2 (.A(in_sample[10]),
    .Y(net2));
 BUFx2_ASAP7_75t_R input1 (.A(in_sample[0]),
    .Y(net1));
 BUFx2_ASAP7_75t_R input13 (.A(in_sample[6]),
    .Y(net13));
 BUFx2_ASAP7_75t_R input14 (.A(in_sample[7]),
    .Y(net14));
 BUFx2_ASAP7_75t_R input15 (.A(in_sample[8]),
    .Y(net15));
 BUFx2_ASAP7_75t_R input16 (.A(in_sample[9]),
    .Y(net16));
 BUFx2_ASAP7_75t_R input17 (.A(in_sample_vld),
    .Y(net17));
 BUFx2_ASAP7_75t_R input18 (.A(out_pred_rdy),
    .Y(net18));
 BUFx16f_ASAP7_75t_R input19 (.A(rst),
    .Y(net19));
 BUFx2_ASAP7_75t_R output20 (.A(net20),
    .Y(in_sample_rdy));
 BUFx2_ASAP7_75t_R output21 (.A(net21),
    .Y(out_pred[0]));
 BUFx2_ASAP7_75t_R output22 (.A(net22),
    .Y(out_pred[10]));
 BUFx2_ASAP7_75t_R output23 (.A(net23),
    .Y(out_pred[11]));
 BUFx2_ASAP7_75t_R output24 (.A(net24),
    .Y(out_pred[12]));
 BUFx2_ASAP7_75t_R output25 (.A(net25),
    .Y(out_pred[13]));
 BUFx2_ASAP7_75t_R output26 (.A(net26),
    .Y(out_pred[14]));
 BUFx2_ASAP7_75t_R output27 (.A(net27),
    .Y(out_pred[15]));
 BUFx2_ASAP7_75t_R output28 (.A(net28),
    .Y(out_pred[1]));
 BUFx2_ASAP7_75t_R output29 (.A(net29),
    .Y(out_pred[2]));
 BUFx2_ASAP7_75t_R output30 (.A(net30),
    .Y(out_pred[3]));
 BUFx2_ASAP7_75t_R output31 (.A(net31),
    .Y(out_pred[4]));
 BUFx2_ASAP7_75t_R output32 (.A(net32),
    .Y(out_pred[5]));
 BUFx2_ASAP7_75t_R output33 (.A(net33),
    .Y(out_pred[6]));
 BUFx2_ASAP7_75t_R output34 (.A(net34),
    .Y(out_pred[7]));
 BUFx2_ASAP7_75t_R output35 (.A(net35),
    .Y(out_pred[8]));
 BUFx2_ASAP7_75t_R output36 (.A(net36),
    .Y(out_pred[9]));
 BUFx2_ASAP7_75t_R output37 (.A(net37),
    .Y(out_pred_vld));
 BUFx16f_ASAP7_75t_R repeater38 (.A(_1507_),
    .Y(net38));
 BUFx16f_ASAP7_75t_R repeater39 (.A(_1507_),
    .Y(net39));
 BUFx12f_ASAP7_75t_R repeater40 (.A(_0820_),
    .Y(net40));
 BUFx10_ASAP7_75t_R repeater41 (.A(net196),
    .Y(net41));
 BUFx10_ASAP7_75t_R repeater42 (.A(net43),
    .Y(net42));
 BUFx10_ASAP7_75t_R repeater43 (.A(_0263_),
    .Y(net43));
 BUFx12f_ASAP7_75t_R repeater44 (.A(_0266_),
    .Y(net44));
 BUFx6f_ASAP7_75t_R repeater45 (.A(_0266_),
    .Y(net45));
 BUFx10_ASAP7_75t_R repeater46 (.A(net210),
    .Y(net46));
 BUFx6f_ASAP7_75t_R repeater47 (.A(net217),
    .Y(net47));
 BUFx10_ASAP7_75t_R repeater48 (.A(_0267_),
    .Y(net48));
 BUFx10_ASAP7_75t_R repeater49 (.A(_0267_),
    .Y(net49));
 INVx2_ASAP7_75t_R _5880__1 (.A(clknet_3_2__leaf_clk),
    .Y(net50));
 INVx2_ASAP7_75t_R _5880__2 (.A(clknet_3_2__leaf_clk),
    .Y(net51));
 INVx2_ASAP7_75t_R _5880__3 (.A(clknet_3_6__leaf_clk),
    .Y(net52));
 INVx2_ASAP7_75t_R _5880__4 (.A(clknet_3_6__leaf_clk),
    .Y(net53));
 INVx2_ASAP7_75t_R _5880__5 (.A(clknet_3_6__leaf_clk),
    .Y(net54));
 INVx2_ASAP7_75t_R _5880__6 (.A(clknet_3_6__leaf_clk),
    .Y(net55));
 INVx2_ASAP7_75t_R _5880__7 (.A(clknet_3_3__leaf_clk),
    .Y(net56));
 INVx2_ASAP7_75t_R _5880__8 (.A(clknet_3_3__leaf_clk),
    .Y(net57));
 INVx2_ASAP7_75t_R _5880__9 (.A(clknet_3_3__leaf_clk),
    .Y(net58));
 INVx2_ASAP7_75t_R _5880__10 (.A(clknet_3_3__leaf_clk),
    .Y(net59));
 INVx2_ASAP7_75t_R _5880__11 (.A(clknet_3_3__leaf_clk),
    .Y(net60));
 INVx2_ASAP7_75t_R _5880__12 (.A(clknet_3_2__leaf_clk),
    .Y(net61));
 INVx2_ASAP7_75t_R _5880__13 (.A(clknet_3_2__leaf_clk),
    .Y(net62));
 INVx2_ASAP7_75t_R _5880__14 (.A(clknet_3_2__leaf_clk),
    .Y(net63));
 INVx2_ASAP7_75t_R _5880__15 (.A(clknet_3_2__leaf_clk),
    .Y(net64));
 INVx2_ASAP7_75t_R _5880__16 (.A(clknet_3_2__leaf_clk),
    .Y(net65));
 INVx2_ASAP7_75t_R _5880__17 (.A(clknet_3_2__leaf_clk),
    .Y(net66));
 INVx2_ASAP7_75t_R _5880__18 (.A(clknet_3_2__leaf_clk),
    .Y(net67));
 INVx2_ASAP7_75t_R _5880__19 (.A(clknet_3_4__leaf_clk),
    .Y(net68));
 INVx2_ASAP7_75t_R _5880__20 (.A(clknet_3_5__leaf_clk),
    .Y(net69));
 INVx2_ASAP7_75t_R _5880__21 (.A(clknet_3_5__leaf_clk),
    .Y(net70));
 INVx2_ASAP7_75t_R _5880__22 (.A(clknet_3_5__leaf_clk),
    .Y(net71));
 INVx2_ASAP7_75t_R _5880__23 (.A(clknet_3_5__leaf_clk),
    .Y(net72));
 INVx2_ASAP7_75t_R _5880__24 (.A(clknet_3_5__leaf_clk),
    .Y(net73));
 INVx2_ASAP7_75t_R _5880__25 (.A(clknet_3_5__leaf_clk),
    .Y(net74));
 INVx2_ASAP7_75t_R _26 (.A(clknet_3_5__leaf_clk),
    .Y(net75));
 INVx2_ASAP7_75t_R _26_27 (.A(clknet_3_5__leaf_clk),
    .Y(net76));
 INVx2_ASAP7_75t_R _26_28 (.A(clknet_3_5__leaf_clk),
    .Y(net77));
 INVx2_ASAP7_75t_R _26_29 (.A(clknet_3_5__leaf_clk),
    .Y(net78));
 INVx2_ASAP7_75t_R _26_30 (.A(clknet_3_5__leaf_clk),
    .Y(net79));
 INVx2_ASAP7_75t_R _26_31 (.A(clknet_3_5__leaf_clk),
    .Y(net80));
 INVx2_ASAP7_75t_R _26_32 (.A(clknet_3_5__leaf_clk),
    .Y(net81));
 INVx2_ASAP7_75t_R _26_33 (.A(clknet_3_5__leaf_clk),
    .Y(net82));
 INVx2_ASAP7_75t_R _26_34 (.A(clknet_3_5__leaf_clk),
    .Y(net83));
 INVx2_ASAP7_75t_R _26_35 (.A(clknet_3_5__leaf_clk),
    .Y(net84));
 INVx2_ASAP7_75t_R _26_36 (.A(clknet_3_4__leaf_clk),
    .Y(net85));
 INVx2_ASAP7_75t_R _26_37 (.A(clknet_3_5__leaf_clk),
    .Y(net86));
 INVx2_ASAP7_75t_R _26_38 (.A(clknet_3_5__leaf_clk),
    .Y(net87));
 INVx2_ASAP7_75t_R _26_39 (.A(clknet_3_4__leaf_clk),
    .Y(net88));
 INVx2_ASAP7_75t_R _26_40 (.A(clknet_3_4__leaf_clk),
    .Y(net89));
 INVx2_ASAP7_75t_R _26_41 (.A(clknet_3_4__leaf_clk),
    .Y(net90));
 INVx2_ASAP7_75t_R _26_42 (.A(clknet_3_4__leaf_clk),
    .Y(net91));
 INVx2_ASAP7_75t_R _26_43 (.A(clknet_3_4__leaf_clk),
    .Y(net92));
 INVx2_ASAP7_75t_R _26_44 (.A(clknet_3_4__leaf_clk),
    .Y(net93));
 INVx2_ASAP7_75t_R _26_45 (.A(clknet_3_4__leaf_clk),
    .Y(net94));
 INVx2_ASAP7_75t_R _26_46 (.A(clknet_3_4__leaf_clk),
    .Y(net95));
 INVx2_ASAP7_75t_R _26_47 (.A(clknet_3_4__leaf_clk),
    .Y(net96));
 INVx2_ASAP7_75t_R _26_48 (.A(clknet_3_4__leaf_clk),
    .Y(net97));
 INVx2_ASAP7_75t_R _26_49 (.A(clknet_3_1__leaf_clk),
    .Y(net98));
 INVx2_ASAP7_75t_R _26_50 (.A(clknet_3_1__leaf_clk),
    .Y(net99));
 INVx2_ASAP7_75t_R _26_51 (.A(clknet_3_1__leaf_clk),
    .Y(net100));
 INVx2_ASAP7_75t_R _26_52 (.A(clknet_3_1__leaf_clk),
    .Y(net101));
 INVx2_ASAP7_75t_R _26_53 (.A(clknet_3_1__leaf_clk),
    .Y(net102));
 INVx2_ASAP7_75t_R _26_54 (.A(clknet_3_1__leaf_clk),
    .Y(net103));
 INVx2_ASAP7_75t_R _26_55 (.A(clknet_3_1__leaf_clk),
    .Y(net104));
 INVx2_ASAP7_75t_R _26_56 (.A(clknet_3_1__leaf_clk),
    .Y(net105));
 INVx2_ASAP7_75t_R _26_57 (.A(clknet_3_1__leaf_clk),
    .Y(net106));
 INVx2_ASAP7_75t_R _26_58 (.A(clknet_3_1__leaf_clk),
    .Y(net107));
 INVx2_ASAP7_75t_R _26_59 (.A(clknet_3_1__leaf_clk),
    .Y(net108));
 INVx2_ASAP7_75t_R _26_60 (.A(clknet_3_0__leaf_clk),
    .Y(net109));
 INVx2_ASAP7_75t_R _26_61 (.A(clknet_3_0__leaf_clk),
    .Y(net110));
 INVx2_ASAP7_75t_R _26_62 (.A(clknet_3_0__leaf_clk),
    .Y(net111));
 INVx2_ASAP7_75t_R _26_63 (.A(clknet_3_0__leaf_clk),
    .Y(net112));
 INVx2_ASAP7_75t_R _26_64 (.A(clknet_3_0__leaf_clk),
    .Y(net113));
 INVx2_ASAP7_75t_R _26_65 (.A(clknet_3_0__leaf_clk),
    .Y(net114));
 INVx2_ASAP7_75t_R _26_66 (.A(clknet_3_0__leaf_clk),
    .Y(net115));
 INVx2_ASAP7_75t_R _26_67 (.A(clknet_3_0__leaf_clk),
    .Y(net116));
 INVx2_ASAP7_75t_R _26_68 (.A(clknet_3_0__leaf_clk),
    .Y(net117));
 INVx2_ASAP7_75t_R _26_69 (.A(clknet_3_0__leaf_clk),
    .Y(net118));
 INVx2_ASAP7_75t_R _26_70 (.A(clknet_3_0__leaf_clk),
    .Y(net119));
 INVx2_ASAP7_75t_R _26_71 (.A(clknet_3_0__leaf_clk),
    .Y(net120));
 INVx2_ASAP7_75t_R _26_72 (.A(clknet_3_0__leaf_clk),
    .Y(net121));
 INVx2_ASAP7_75t_R _26_73 (.A(clknet_3_0__leaf_clk),
    .Y(net122));
 INVx2_ASAP7_75t_R _26_74 (.A(clknet_3_0__leaf_clk),
    .Y(net123));
 INVx2_ASAP7_75t_R _26_75 (.A(clknet_3_0__leaf_clk),
    .Y(net124));
 INVx2_ASAP7_75t_R _76 (.A(clknet_3_0__leaf_clk),
    .Y(net125));
 INVx2_ASAP7_75t_R _76_77 (.A(clknet_3_0__leaf_clk),
    .Y(net126));
 INVx2_ASAP7_75t_R _76_78 (.A(clknet_3_1__leaf_clk),
    .Y(net127));
 INVx2_ASAP7_75t_R _76_79 (.A(clknet_3_0__leaf_clk),
    .Y(net128));
 INVx2_ASAP7_75t_R _76_80 (.A(clknet_3_1__leaf_clk),
    .Y(net129));
 INVx2_ASAP7_75t_R _76_81 (.A(clknet_3_7__leaf_clk),
    .Y(net130));
 INVx2_ASAP7_75t_R _76_82 (.A(clknet_3_7__leaf_clk),
    .Y(net131));
 INVx2_ASAP7_75t_R _76_83 (.A(clknet_3_7__leaf_clk),
    .Y(net132));
 INVx2_ASAP7_75t_R _76_84 (.A(clknet_3_7__leaf_clk),
    .Y(net133));
 INVx2_ASAP7_75t_R _76_85 (.A(clknet_3_7__leaf_clk),
    .Y(net134));
 INVx2_ASAP7_75t_R _76_86 (.A(clknet_3_7__leaf_clk),
    .Y(net135));
 INVx2_ASAP7_75t_R _76_87 (.A(clknet_3_7__leaf_clk),
    .Y(net136));
 INVx2_ASAP7_75t_R _76_88 (.A(clknet_3_7__leaf_clk),
    .Y(net137));
 INVx2_ASAP7_75t_R _76_89 (.A(clknet_3_7__leaf_clk),
    .Y(net138));
 INVx2_ASAP7_75t_R _76_90 (.A(clknet_3_7__leaf_clk),
    .Y(net139));
 INVx2_ASAP7_75t_R _76_91 (.A(clknet_3_7__leaf_clk),
    .Y(net140));
 INVx2_ASAP7_75t_R _76_92 (.A(clknet_3_7__leaf_clk),
    .Y(net141));
 INVx2_ASAP7_75t_R _76_93 (.A(clknet_3_7__leaf_clk),
    .Y(net142));
 INVx2_ASAP7_75t_R _76_94 (.A(clknet_3_7__leaf_clk),
    .Y(net143));
 INVx2_ASAP7_75t_R _76_95 (.A(clknet_3_7__leaf_clk),
    .Y(net144));
 INVx2_ASAP7_75t_R _76_96 (.A(clknet_3_6__leaf_clk),
    .Y(net145));
 INVx2_ASAP7_75t_R _76_97 (.A(clknet_3_6__leaf_clk),
    .Y(net146));
 INVx2_ASAP7_75t_R _76_98 (.A(clknet_3_6__leaf_clk),
    .Y(net147));
 INVx2_ASAP7_75t_R _76_99 (.A(clknet_3_6__leaf_clk),
    .Y(net148));
 INVx2_ASAP7_75t_R _76_100 (.A(clknet_3_6__leaf_clk),
    .Y(net149));
 INVx2_ASAP7_75t_R _76_101 (.A(clknet_3_6__leaf_clk),
    .Y(net150));
 INVx2_ASAP7_75t_R _76_102 (.A(clknet_3_3__leaf_clk),
    .Y(net151));
 INVx2_ASAP7_75t_R _76_103 (.A(clknet_3_3__leaf_clk),
    .Y(net152));
 INVx2_ASAP7_75t_R _76_104 (.A(clknet_3_3__leaf_clk),
    .Y(net153));
 INVx2_ASAP7_75t_R _76_105 (.A(clknet_3_3__leaf_clk),
    .Y(net154));
 INVx2_ASAP7_75t_R _76_106 (.A(clknet_3_3__leaf_clk),
    .Y(net155));
 INVx2_ASAP7_75t_R _76_107 (.A(clknet_3_3__leaf_clk),
    .Y(net156));
 INVx2_ASAP7_75t_R _76_108 (.A(clknet_3_2__leaf_clk),
    .Y(net157));
 INVx2_ASAP7_75t_R _76_109 (.A(clknet_3_2__leaf_clk),
    .Y(net158));
 INVx2_ASAP7_75t_R _76_110 (.A(clknet_3_2__leaf_clk),
    .Y(net159));
 INVx2_ASAP7_75t_R _76_111 (.A(clknet_3_2__leaf_clk),
    .Y(net160));
 INVx2_ASAP7_75t_R _76_112 (.A(clknet_3_2__leaf_clk),
    .Y(net161));
 BUFx4_ASAP7_75t_R clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .Y(clknet_3_0__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .Y(clknet_3_1__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .Y(clknet_3_2__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .Y(clknet_3_3__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .Y(clknet_3_4__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .Y(clknet_3_5__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .Y(clknet_3_6__leaf_clk));
 BUFx4_ASAP7_75t_R clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .Y(clknet_3_7__leaf_clk));
 BUFx16f_ASAP7_75t_R split113 (.A(net195),
    .Y(net162));
 BUFx3_ASAP7_75t_R rebuffer114 (.A(_0714_),
    .Y(net163));
 BUFx2_ASAP7_75t_R rebuffer115 (.A(net163),
    .Y(net164));
 BUFx2_ASAP7_75t_R rebuffer116 (.A(net163),
    .Y(net165));
 BUFx2_ASAP7_75t_R rebuffer117 (.A(net163),
    .Y(net166));
 BUFx2_ASAP7_75t_R rebuffer118 (.A(net163),
    .Y(net167));
 BUFx2_ASAP7_75t_R rebuffer119 (.A(net167),
    .Y(net168));
 BUFx3_ASAP7_75t_R rebuffer120 (.A(_0025_),
    .Y(net169));
 BUFx2_ASAP7_75t_R rebuffer121 (.A(net169),
    .Y(net170));
 BUFx2_ASAP7_75t_R rebuffer122 (.A(net169),
    .Y(net171));
 BUFx2_ASAP7_75t_R rebuffer123 (.A(net169),
    .Y(net172));
 BUFx2_ASAP7_75t_R rebuffer124 (.A(_0430_),
    .Y(net173));
 BUFx2_ASAP7_75t_R rebuffer125 (.A(_0430_),
    .Y(net174));
 BUFx2_ASAP7_75t_R rebuffer126 (.A(net174),
    .Y(net175));
 BUFx3_ASAP7_75t_R rebuffer127 (.A(_0710_),
    .Y(net176));
 BUFx2_ASAP7_75t_R rebuffer128 (.A(net176),
    .Y(net177));
 BUFx2_ASAP7_75t_R rebuffer129 (.A(net176),
    .Y(net178));
 BUFx2_ASAP7_75t_R rebuffer130 (.A(net176),
    .Y(net179));
 BUFx16f_ASAP7_75t_R split131 (.A(net209),
    .Y(net180));
 BUFx3_ASAP7_75t_R rebuffer132 (.A(_0711_),
    .Y(net181));
 BUFx2_ASAP7_75t_R rebuffer133 (.A(net181),
    .Y(net182));
 BUFx2_ASAP7_75t_R rebuffer134 (.A(net182),
    .Y(net183));
 BUFx2_ASAP7_75t_R rebuffer135 (.A(net181),
    .Y(net184));
 BUFx2_ASAP7_75t_R rebuffer136 (.A(net181),
    .Y(net185));
 BUFx2_ASAP7_75t_R rebuffer137 (.A(_0743_),
    .Y(net186));
 BUFx2_ASAP7_75t_R rebuffer138 (.A(_0743_),
    .Y(net187));
 BUFx2_ASAP7_75t_R rebuffer139 (.A(net187),
    .Y(net188));
 BUFx2_ASAP7_75t_R rebuffer140 (.A(net188),
    .Y(net189));
 BUFx3_ASAP7_75t_R rebuffer141 (.A(_0715_),
    .Y(net190));
 BUFx2_ASAP7_75t_R rebuffer142 (.A(net190),
    .Y(net191));
 BUFx2_ASAP7_75t_R rebuffer143 (.A(net191),
    .Y(net192));
 BUFx2_ASAP7_75t_R rebuffer144 (.A(net190),
    .Y(net193));
 BUFx2_ASAP7_75t_R rebuffer145 (.A(net190),
    .Y(net194));
 BUFx12_ASAP7_75t_R split146 (.A(net227),
    .Y(net195));
 BUFx3_ASAP7_75t_R rebuffer147 (.A(_0699_),
    .Y(net196));
 BUFx2_ASAP7_75t_R rebuffer148 (.A(net196),
    .Y(net197));
 BUFx2_ASAP7_75t_R rebuffer149 (.A(net196),
    .Y(net198));
 BUFx2_ASAP7_75t_R rebuffer150 (.A(net196),
    .Y(net199));
 BUFx2_ASAP7_75t_R rebuffer151 (.A(net199),
    .Y(net200));
 BUFx2_ASAP7_75t_R rebuffer152 (.A(net196),
    .Y(net201));
 BUFx6f_ASAP7_75t_R rebuffer153 (.A(net201),
    .Y(net202));
 BUFx2_ASAP7_75t_R rebuffer154 (.A(net202),
    .Y(net203));
 BUFx2_ASAP7_75t_R rebuffer155 (.A(net202),
    .Y(net204));
 BUFx2_ASAP7_75t_R rebuffer156 (.A(net204),
    .Y(net205));
 BUFx3_ASAP7_75t_R rebuffer157 (.A(_0716_),
    .Y(net206));
 BUFx2_ASAP7_75t_R rebuffer158 (.A(net206),
    .Y(net207));
 BUFx2_ASAP7_75t_R rebuffer159 (.A(net206),
    .Y(net208));
 BUFx10_ASAP7_75t_R split160 (.A(_1173_),
    .Y(net209));
 BUFx3_ASAP7_75t_R rebuffer161 (.A(_0696_),
    .Y(net210));
 BUFx2_ASAP7_75t_R rebuffer162 (.A(net210),
    .Y(net211));
 BUFx6f_ASAP7_75t_R rebuffer163 (.A(net211),
    .Y(net212));
 BUFx2_ASAP7_75t_R rebuffer164 (.A(net212),
    .Y(net213));
 BUFx2_ASAP7_75t_R rebuffer165 (.A(net212),
    .Y(net214));
 BUFx2_ASAP7_75t_R rebuffer166 (.A(net212),
    .Y(net215));
 BUFx2_ASAP7_75t_R rebuffer167 (.A(net210),
    .Y(net216));
 BUFx2_ASAP7_75t_R rebuffer168 (.A(net210),
    .Y(net217));
 BUFx2_ASAP7_75t_R rebuffer169 (.A(net210),
    .Y(net218));
 BUFx12_ASAP7_75t_R split170 (.A(net221),
    .Y(net219));
 BUFx2_ASAP7_75t_R rebuffer171 (.A(_0744_),
    .Y(net220));
 BUFx6f_ASAP7_75t_R split172 (.A(_1676_),
    .Y(net221));
 BUFx16f_ASAP7_75t_R split173 (.A(net228),
    .Y(net222));
 BUFx6f_ASAP7_75t_R split174 (.A(net233),
    .Y(net223));
 BUFx4f_ASAP7_75t_R split175 (.A(_2871_),
    .Y(net224));
 BUFx2_ASAP7_75t_R split176 (.A(_1676_),
    .Y(net225));
 BUFx6f_ASAP7_75t_R split177 (.A(net234),
    .Y(net226));
 BUFx6f_ASAP7_75t_R split178 (.A(net237),
    .Y(net227));
 BUFx10_ASAP7_75t_R split179 (.A(net236),
    .Y(net228));
 BUFx16f_ASAP7_75t_R split180 (.A(_1508_),
    .Y(net229));
 BUFx2_ASAP7_75t_R rebuffer181 (.A(_0745_),
    .Y(net230));
 BUFx2_ASAP7_75t_R rebuffer182 (.A(net230),
    .Y(net231));
 BUFx2_ASAP7_75t_R rebuffer183 (.A(net231),
    .Y(net232));
 BUFx3_ASAP7_75t_R split184 (.A(_1507_),
    .Y(net233));
 BUFx3_ASAP7_75t_R split185 (.A(_1674_),
    .Y(net234));
 BUFx6f_ASAP7_75t_R rebuffer186 (.A(_2871_),
    .Y(net235));
 BUFx4f_ASAP7_75t_R split187 (.A(_1864_),
    .Y(net236));
 BUFx3_ASAP7_75t_R split188 (.A(_1178_),
    .Y(net237));
 BUFx2_ASAP7_75t_R rebuffer189 (.A(_0452_),
    .Y(net238));
 BUFx2_ASAP7_75t_R rebuffer190 (.A(_1178_),
    .Y(net239));
 FILLERxp5_ASAP7_75t_R FILLER_0_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_75 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_76 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_77 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_64 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_67 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_92 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_3 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_5 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_28 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_31 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_35 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_36 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_37 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_38 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_41 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_42 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_43 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_44 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_47 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_49 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_50 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_52 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_55 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_69 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_70 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_83 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_84 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_86 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_212 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_515 ();
endmodule
